module patch (t_0, t_1, t_2, t_3, t_4, t_5, t_6, t_7, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13;
output t_0, t_1, t_2, t_3, t_4, t_5, t_6, t_7;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238;

nor ( w1 , g3 , g4 );
nor ( w2 , g6 , g7 );
and ( w3 , g5 , w6535 );
and ( w4 , w1 , w3 );
and ( w5 , w7102 , g3 );
and ( w6 , g5 , g6 );
and ( w7 , g7 , g5 );
nor ( w8 , w6 , w7 );
nor ( w9 , w8 , w3 );
nor ( w10 , w5 , w9 );
and ( w11 , g6 , w7104 );
nor ( w12 , g7 , w11 );
nor ( w13 , w12 , w8 );
and ( w14 , w10 , w1025 );
nor ( w15 , g8 , g9 );
nor ( w16 , w14 , w15 );
not ( w17 , w4 );
and ( w18 , w17 , w16 );
and ( w19 , w5 , w403 );
and ( w20 , w19 , w1025 );
nor ( w21 , w20 , g10 );
not ( w22 , w21 );
and ( w23 , w22 , g2 );
nor ( w24 , w23 , g10 );
and ( w25 , w18 , w24 );
and ( w26 , w25 , w6945 );
and ( w27 , w3 , g3 );
and ( w28 , w3 , w7097 );
nor ( w29 , w28 , w15 );
not ( w30 , w27 );
and ( w31 , w30 , w29 );
not ( w32 , w31 );
and ( w33 , w32 , g4 );
not ( w34 , w20 );
and ( w35 , w34 , g1 );
and ( w36 , w35 , w6997 );
not ( w37 , w33 );
and ( w38 , w37 , w36 );
and ( w39 , w38 , w7183 );
nor ( w40 , w26 , w39 );
and ( w41 , w40 , g2 );
nor ( w42 , w9 , w13 );
not ( w43 , w42 );
and ( w44 , w43 , g1 );
and ( w45 , w44 , w6997 );
and ( w46 , w4497 , g4 );
and ( w47 , g1 , w6794 );
and ( w48 , w47 , w7183 );
and ( w49 , w48 , w6997 );
nor ( w50 , w49 , g4 );
nor ( w51 , w50 , w15 );
and ( w52 , w51 , w6997 );
not ( w53 , w46 );
and ( w54 , w53 , w52 );
not ( w55 , w54 );
and ( w56 , w55 , g3 );
and ( w57 , g1 , g4 );
and ( w58 , w57 , w6794 );
and ( w59 , w58 , w7183 );
and ( w60 , w59 , w6997 );
nor ( w61 , w44 , w60 );
and ( w62 , w7102 , w3 );
nor ( w63 , w62 , w15 );
not ( w64 , w61 );
and ( w65 , w64 , w63 );
nor ( w66 , w65 , g3 );
and ( w67 , w66 , w7213 );
nor ( w68 , w67 , w15 );
and ( w69 , w68 , w6997 );
not ( w70 , w56 );
and ( w71 , w70 , w69 );
nor ( w72 , w71 , g2 );
nor ( w73 , w72 , w15 );
and ( w74 , w73 , w6997 );
not ( w75 , w41 );
and ( w76 , w75 , w74 );
and ( w77 , w76 , w7094 );
and ( w78 , w6380 , g1 );
and ( w79 , g1 , w6471 );
nor ( w80 , w79 , w13 );
not ( w81 , w80 );
and ( w82 , w81 , g12 );
and ( w83 , w82 , g1 );
nor ( w84 , w78 , w83 );
nor ( w85 , w84 , g3 );
and ( w86 , w85 , g11 );
nor ( w87 , g7 , w8 );
nor ( w88 , w87 , w9 );
nor ( w89 , w88 , g6 );
nor ( w90 , g2 , w89 );
not ( w91 , w90 );
and ( w92 , w91 , g4 );
and ( w93 , w92 , w7183 );
and ( w94 , g2 , g3 );
and ( w95 , w6471 , g4 );
and ( w96 , w95 , w15 );
and ( w97 , w96 , g1 );
and ( w98 , w97 , w6997 );
and ( w99 , w98 , w6794 );
nor ( w100 , w99 , w13 );
nor ( w101 , w100 , g3 );
and ( w102 , w101 , w7213 );
and ( w103 , w102 , w15 );
nor ( w104 , w103 , g10 );
not ( w105 , w104 );
and ( w106 , w105 , g11 );
nor ( w107 , w106 , g2 );
nor ( w108 , w107 , g3 );
and ( w109 , w108 , w15 );
and ( w110 , w109 , w6471 );
and ( w111 , w110 , g11 );
nor ( w112 , w94 , w111 );
nor ( w113 , w112 , w3 );
and ( w114 , w113 , g4 );
and ( w115 , w114 , w15 );
and ( w116 , w115 , w6471 );
nor ( w117 , w116 , g10 );
not ( w118 , w117 );
and ( w119 , w118 , g11 );
nor ( w120 , w119 , g10 );
and ( w121 , w4009 , w120 );
and ( w122 , w121 , w3 );
and ( w123 , g1 , g11 );
not ( w124 , w123 );
and ( w125 , g11 , w124 );
and ( w126 , w125 , g13 );
and ( w127 , w126 , g4 );
and ( w128 , w127 , g2 );
and ( w129 , g11 , w99 );
and ( w130 , w129 , w7213 );
and ( w131 , w130 , w7097 );
not ( w132 , w131 );
and ( w133 , g11 , w132 );
not ( w134 , w133 );
and ( w135 , w134 , g4 );
and ( w136 , w135 , w7213 );
and ( w137 , w136 , w6997 );
and ( w138 , w137 , w7097 );
and ( w139 , w138 , w6794 );
nor ( w140 , w128 , w139 );
nor ( w141 , w140 , g10 );
and ( w142 , w141 , w7097 );
and ( w143 , w142 , w15 );
and ( w144 , w143 , w6794 );
and ( w145 , w144 , g11 );
and ( w146 , w111 , g4 );
and ( w147 , g1 , w7213 );
and ( w148 , w6997 , g2 );
and ( w149 , w15 , w403 );
and ( w150 , w149 , w1025 );
and ( w151 , w7213 , w150 );
and ( w152 , w151 , w7102 );
and ( w153 , w152 , g3 );
nor ( w154 , w148 , w153 );
nor ( w155 , w154 , g4 );
and ( w156 , w155 , w1025 );
and ( w157 , w156 , g3 );
and ( w158 , w147 , w848 );
and ( w159 , w158 , g3 );
and ( w160 , g1 , g2 );
and ( w161 , w160 , w7097 );
and ( w162 , w161 , w7183 );
not ( w163 , w162 );
and ( w164 , w163 , w8 );
nor ( w165 , w164 , w3 );
nor ( w166 , w165 , g10 );
nor ( w167 , w166 , g4 );
and ( w168 , w167 , g11 );
nor ( w169 , w159 , w168 );
and ( w170 , w169 , g12 );
nor ( w171 , w170 , w15 );
and ( w172 , g4 , w7183 );
and ( w173 , w172 , w6794 );
and ( w174 , w173 , g10 );
and ( w175 , g3 , g4 );
and ( w176 , w175 , w6794 );
and ( w177 , w176 , w15 );
and ( w178 , w177 , g10 );
nor ( w179 , w174 , w178 );
and ( w180 , w179 , g2 );
nor ( w181 , g3 , w180 );
and ( w182 , w5 , w7183 );
nor ( w183 , w181 , w182 );
nor ( w184 , w183 , w3 );
and ( w185 , w184 , g10 );
nor ( w186 , w185 , w178 );
and ( w187 , w186 , g2 );
not ( w188 , w187 );
and ( w189 , w188 , g10 );
and ( w190 , w1 , w6997 );
nor ( w191 , w190 , w178 );
and ( w192 , w191 , g2 );
not ( w193 , w175 );
and ( w194 , w193 , w192 );
nor ( w195 , w194 , w3 );
and ( w196 , w195 , w6997 );
not ( w197 , w196 );
and ( w198 , w197 , g2 );
and ( w199 , w198 , g11 );
nor ( w200 , w199 , w15 );
and ( w201 , w175 , w3795 );
and ( w202 , w3555 , g2 );
and ( w203 , w536 , w202 );
not ( w204 , w203 );
and ( w205 , w204 , w15 );
and ( w206 , w205 , w6997 );
not ( w207 , w206 );
and ( w208 , w207 , g2 );
and ( w209 , w208 , g11 );
not ( w210 , w200 );
and ( w211 , w210 , w209 );
and ( w212 , w211 , w470 );
not ( w213 , w189 );
and ( w214 , w213 , w212 );
nor ( w215 , w3 , w15 );
and ( w216 , w1025 , w3 );
and ( w217 , w475 , w15 );
nor ( w218 , w215 , w217 );
nor ( w219 , w218 , g10 );
nor ( w220 , w219 , g2 );
and ( w221 , w215 , g10 );
not ( w222 , w221 );
and ( w223 , w220 , w222 );
not ( w224 , w223 );
and ( w225 , w224 , g3 );
nor ( w226 , g10 , w9 );
nor ( w227 , w226 , w15 );
nor ( w228 , w7 , w11 );
nor ( w229 , w228 , g13 );
and ( w230 , g13 , g1 );
nor ( w231 , g13 , g1 );
nor ( w232 , w230 , w231 );
nor ( w233 , w232 , w8 );
and ( w234 , g13 , w6794 );
and ( w235 , w6945 , w234 );
and ( w236 , w235 , g10 );
nor ( w237 , w233 , w236 );
not ( w238 , w237 );
and ( w239 , w238 , g10 );
and ( w240 , g1 , w6997 );
and ( w241 , w6997 , w13 );
and ( w242 , g10 , w6945 );
nor ( w243 , w7 , g13 );
and ( w244 , w243 , g1 );
and ( w245 , w244 , w6997 );
and ( w246 , w245 , w5796 );
and ( w247 , w246 , w5798 );
nor ( w248 , w242 , w247 );
nor ( w249 , w248 , g13 );
and ( w250 , w249 , w5796 );
and ( w251 , w250 , w5798 );
nor ( w252 , w241 , w251 );
nor ( w253 , w45 , w245 );
and ( w254 , w253 , w7102 );
nor ( w255 , w254 , g8 );
and ( w256 , w255 , w5798 );
not ( w257 , w252 );
and ( w258 , w257 , w256 );
nor ( w259 , w240 , w258 );
nor ( w260 , w259 , g10 );
and ( w261 , w260 , w15 );
nor ( w262 , w239 , w261 );
not ( w263 , w262 );
and ( w264 , w263 , w15 );
nor ( w265 , w229 , w264 );
not ( w266 , w265 );
and ( w267 , w266 , w15 );
and ( w268 , w267 , w7097 );
and ( w269 , w268 , w7213 );
and ( w270 , w269 , g10 );
not ( w271 , w270 );
and ( w272 , w271 , w3 );
nor ( w273 , w272 , w8 );
not ( w274 , w273 );
and ( w275 , w274 , g11 );
not ( w276 , w227 );
and ( w277 , w276 , w275 );
and ( w278 , w277 , w3 );
and ( w279 , w12 , g5 );
nor ( w280 , w279 , w8 );
not ( w281 , w278 );
and ( w282 , w281 , w280 );
and ( w283 , w240 , w15 );
and ( w284 , w283 , w6794 );
not ( w285 , w284 );
and ( w286 , w285 , g11 );
not ( w287 , w282 );
and ( w288 , w287 , w286 );
nor ( w289 , w288 , g3 );
nor ( w290 , w289 , w144 );
and ( w291 , w290 , w7213 );
and ( w292 , w291 , g11 );
not ( w293 , w225 );
and ( w294 , w293 , w292 );
and ( w295 , w294 , g4 );
and ( w296 , g10 , w13 );
nor ( w297 , w296 , w9 );
not ( w298 , w297 );
and ( w299 , w298 , g3 );
and ( w300 , w299 , w7183 );
nor ( w301 , w216 , g3 );
and ( w302 , w301 , g10 );
and ( w303 , w302 , w13 );
and ( w304 , g10 , g3 );
and ( w305 , w304 , w6794 );
and ( w306 , w305 , w15 );
nor ( w307 , w303 , w306 );
not ( w308 , w307 );
and ( w309 , w308 , w15 );
nor ( w310 , w300 , w309 );
and ( w311 , w42 , g3 );
and ( w312 , w311 , w6997 );
and ( w313 , w312 , w7183 );
and ( w314 , g3 , w6997 );
and ( w315 , w314 , w280 );
and ( w316 , w315 , w15 );
nor ( w317 , w313 , w316 );
and ( w318 , w310 , w317 );
and ( w319 , w318 , w536 );
and ( w320 , w319 , w7102 );
and ( w321 , w320 , w7213 );
nor ( w322 , w295 , w321 );
and ( w323 , w94 , w7102 );
nor ( w324 , w323 , w15 );
nor ( w325 , w280 , w9 );
not ( w326 , w325 );
and ( w327 , w326 , g10 );
and ( w328 , w94 , w15 );
nor ( w329 , w328 , g10 );
nor ( w330 , w327 , w329 );
and ( w331 , w330 , g3 );
and ( w332 , w331 , w15 );
and ( w333 , w332 , w7102 );
and ( w334 , g10 , g4 );
nor ( w335 , w333 , w334 );
and ( w336 , w335 , g2 );
not ( w337 , w336 );
and ( w338 , w337 , g3 );
not ( w339 , w269 );
and ( w340 , w339 , g10 );
not ( w341 , w340 );
and ( w342 , w341 , w15 );
not ( w343 , w342 );
and ( w344 , w343 , w3 );
not ( w345 , w344 );
and ( w346 , w345 , w280 );
not ( w347 , w346 );
and ( w348 , w347 , g10 );
nor ( w349 , w348 , g2 );
and ( w350 , w349 , w15 );
and ( w351 , w350 , w280 );
not ( w352 , w351 );
and ( w353 , w338 , w352 );
nor ( w354 , w329 , g4 );
and ( w355 , w354 , w7097 );
not ( w356 , w355 );
and ( w357 , w356 , g2 );
nor ( w358 , w357 , w351 );
not ( w359 , w358 );
and ( w360 , w359 , w15 );
and ( w361 , w360 , w280 );
not ( w362 , w353 );
and ( w363 , w362 , w361 );
nor ( w364 , w324 , w363 );
not ( w365 , w364 );
and ( w366 , w365 , w280 );
nor ( w367 , g3 , g2 );
and ( w368 , w367 , g10 );
and ( w369 , w368 , w7183 );
and ( w370 , g3 , w7213 );
and ( w371 , w370 , w15 );
not ( w372 , w371 );
and ( w373 , w372 , g4 );
and ( w374 , g10 , w15 );
nor ( w375 , w374 , w332 );
and ( w376 , w375 , g2 );
and ( w377 , w314 , w15 );
nor ( w378 , w377 , g2 );
and ( w379 , w378 , w6794 );
nor ( w380 , w376 , w379 );
nor ( w381 , w380 , w3 );
nor ( w382 , w373 , w381 );
nor ( w383 , w382 , w3 );
not ( w384 , w369 );
and ( w385 , w384 , w383 );
nor ( w386 , w366 , w385 );
and ( w387 , w386 , g11 );
not ( w388 , w387 );
and ( w389 , w322 , w388 );
not ( w390 , w389 );
and ( w391 , w390 , g11 );
nor ( w392 , w214 , w391 );
and ( w393 , w392 , w7097 );
not ( w394 , w393 );
and ( w395 , w394 , g11 );
not ( w396 , w395 );
and ( w397 , g1 , w396 );
and ( w398 , w397 , g11 );
nor ( w399 , w159 , w398 );
nor ( w400 , w399 , w15 );
and ( w401 , w7213 , w15 );
and ( w402 , w4304 , w157 );
not ( w403 , w9 );
and ( w404 , w402 , w403 );
and ( w405 , w404 , w6471 );
not ( w406 , w405 );
and ( w407 , w406 , g3 );
and ( w408 , w146 , w6794 );
nor ( w409 , w408 , g10 );
not ( w410 , w47 );
and ( w411 , w410 , w409 );
nor ( w412 , w411 , g3 );
and ( w413 , w412 , w15 );
not ( w414 , w413 );
and ( w415 , w414 , g12 );
nor ( w416 , w415 , g13 );
and ( w417 , w416 , w7102 );
nor ( w418 , w417 , g10 );
not ( w419 , w418 );
and ( w420 , w419 , g11 );
nor ( w421 , w407 , w420 );
not ( w422 , w421 );
and ( w423 , w422 , w15 );
and ( w424 , w423 , w6471 );
and ( w425 , w424 , w7102 );
and ( w426 , w425 , w6794 );
and ( w427 , w426 , g11 );
nor ( w428 , w400 , w427 );
and ( w429 , w428 , g12 );
nor ( w430 , w429 , g13 );
and ( w431 , w430 , w7102 );
not ( w432 , w431 );
and ( w433 , w432 , w8 );
nor ( w434 , w433 , w3 );
nor ( w435 , w434 , g10 );
not ( w436 , w435 );
and ( w437 , w436 , g11 );
nor ( w438 , w171 , w437 );
nor ( w439 , w438 , g13 );
not ( w440 , w439 );
and ( w441 , w440 , w8 );
nor ( w442 , w441 , w3 );
nor ( w443 , w442 , g10 );
nor ( w444 , w443 , g4 );
and ( w445 , w444 , g11 );
nor ( w446 , w146 , w445 );
and ( w447 , w446 , w1025 );
and ( w448 , w447 , w6997 );
and ( w449 , w1004 , w448 );
nor ( w450 , w122 , w449 );
nor ( w451 , w450 , g1 );
nor ( w452 , w15 , g4 );
nor ( w453 , w452 , g3 );
nor ( w454 , w453 , w15 );
and ( w455 , w454 , w7102 );
and ( w456 , w455 , w470 );
and ( w457 , w456 , g2 );
and ( w458 , w457 , g11 );
nor ( w459 , w458 , w387 );
not ( w460 , w459 );
and ( w461 , w460 , w3 );
not ( w462 , w461 );
and ( w463 , w462 , w280 );
nor ( w464 , w463 , w392 );
not ( w465 , w464 );
and ( w466 , w465 , g10 );
nor ( w467 , w212 , w391 );
and ( w468 , w467 , w6997 );
nor ( w469 , w466 , w468 );
not ( w470 , w178 );
and ( w471 , w469 , w470 );
and ( w472 , w471 , g2 );
nor ( w473 , w472 , w391 );
and ( w474 , w956 , g1 );
not ( w475 , w216 );
and ( w476 , w475 , g4 );
and ( w477 , w476 , w6794 );
nor ( w478 , w477 , w13 );
and ( w479 , w7183 , w478 );
and ( w480 , w479 , w6997 );
nor ( w481 , w480 , g3 );
and ( w482 , w481 , g11 );
nor ( w483 , w15 , w482 );
and ( w484 , w7102 , g2 );
and ( w485 , w484 , w3 );
and ( w486 , w477 , w15 );
and ( w487 , w486 , w6997 );
nor ( w488 , w485 , w487 );
not ( w489 , w488 );
and ( w490 , w489 , w15 );
and ( w491 , w490 , w6997 );
nor ( w492 , w483 , w491 );
and ( w493 , w7102 , w15 );
and ( w494 , w493 , g2 );
not ( w495 , w494 );
and ( w496 , w495 , w13 );
and ( w497 , w15 , w1023 );
not ( w498 , w497 );
and ( w499 , w498 , g4 );
and ( w500 , w499 , w6794 );
nor ( w501 , w500 , w445 );
nor ( w502 , w501 , g3 );
and ( w503 , w502 , g11 );
nor ( w504 , w496 , w503 );
and ( w505 , w504 , w6471 );
and ( w506 , w505 , w6997 );
nor ( w507 , w506 , g3 );
and ( w508 , w507 , g11 );
and ( w509 , w492 , w508 );
not ( w510 , w509 );
and ( w511 , w510 , g12 );
nor ( w512 , w511 , g3 );
and ( w513 , w512 , g11 );
not ( w514 , w513 );
and ( w515 , w474 , w514 );
and ( w516 , w515 , w6997 );
not ( w517 , w516 );
and ( w518 , w517 , g11 );
not ( w519 , w451 );
and ( w520 , w519 , w518 );
not ( w521 , w520 );
and ( w522 , w521 , g12 );
and ( w523 , w522 , w6997 );
nor ( w524 , w523 , g3 );
and ( w525 , w524 , g11 );
nor ( w526 , w15 , g1 );
and ( w527 , w7183 , g13 );
and ( w528 , w6194 , g1 );
and ( w529 , w528 , w280 );
and ( w530 , w529 , w6997 );
and ( w531 , w530 , g11 );
nor ( w532 , w526 , w531 );
and ( w533 , w532 , w3 );
not ( w534 , w533 );
and ( w535 , w534 , w280 );
not ( w536 , w144 );
and ( w537 , g13 , w536 );
not ( w538 , w537 );
and ( w539 , w538 , w15 );
and ( w540 , w539 , w6794 );
and ( w541 , w15 , w956 );
not ( w542 , w541 );
and ( w543 , w542 , g1 );
nor ( w544 , w540 , w543 );
nor ( w545 , w544 , w3 );
and ( w546 , w545 , g2 );
and ( w547 , w546 , w6997 );
nor ( w548 , w547 , g12 );
not ( w549 , w548 );
and ( w550 , w549 , g11 );
nor ( w551 , w535 , w550 );
not ( w552 , w551 );
and ( w553 , w552 , g2 );
and ( w554 , w6945 , g4 );
and ( w555 , g1 , w7102 );
and ( w556 , w555 , g11 );
nor ( w557 , w554 , w556 );
not ( w558 , w557 );
and ( w559 , w558 , w15 );
nor ( w560 , w559 , g12 );
not ( w561 , w560 );
and ( w562 , w561 , g11 );
nor ( w563 , w57 , w562 );
nor ( w564 , w563 , w8 );
and ( w565 , g1 , w7183 );
nor ( w566 , g1 , w139 );
not ( w567 , w566 );
and ( w568 , w567 , w15 );
not ( w569 , w568 );
and ( w570 , w569 , w8 );
nor ( w571 , w570 , w3 );
and ( w572 , w571 , w7213 );
nor ( w573 , w572 , g10 );
nor ( w574 , w573 , g3 );
nor ( w575 , w565 , w574 );
not ( w576 , w575 );
and ( w577 , w576 , g4 );
nor ( w578 , g1 , g12 );
nor ( w579 , w578 , g13 );
and ( w580 , w579 , w437 );
and ( w581 , w580 , w7102 );
and ( w582 , w581 , w6794 );
nor ( w583 , w582 , g10 );
not ( w584 , w583 );
and ( w585 , w584 , g11 );
nor ( w586 , g13 , w585 );
and ( w587 , w586 , w7102 );
not ( w588 , w587 );
and ( w589 , w588 , g11 );
and ( w590 , w7102 , w589 );
not ( w591 , w590 );
and ( w592 , w15 , w591 );
and ( w593 , w592 , w6997 );
not ( w594 , w593 );
and ( w595 , g1 , w594 );
and ( w596 , w595 , w15 );
nor ( w597 , w596 , g10 );
and ( w598 , w597 , g13 );
and ( w599 , w4437 , w445 );
nor ( w600 , w599 , g13 );
and ( w601 , w600 , w6997 );
nor ( w602 , w601 , g3 );
and ( w603 , w602 , g11 );
not ( w604 , w598 );
and ( w605 , w604 , w603 );
and ( w606 , w605 , w7102 );
not ( w607 , w606 );
and ( w608 , w607 , w8 );
nor ( w609 , w608 , w3 );
nor ( w610 , w609 , g12 );
and ( w611 , w610 , w6997 );
nor ( w612 , w611 , g3 );
nor ( w613 , w577 , w612 );
and ( w614 , w613 , w8 );
nor ( w615 , w614 , w3 );
and ( w616 , w615 , w7213 );
nor ( w617 , w616 , g12 );
and ( w618 , w617 , w6997 );
nor ( w619 , w618 , g3 );
and ( w620 , w619 , g11 );
nor ( w621 , w564 , w620 );
nor ( w622 , w621 , g2 );
nor ( w623 , w622 , g12 );
and ( w624 , w623 , w6997 );
nor ( w625 , w624 , g3 );
and ( w626 , w625 , g11 );
nor ( w627 , w553 , w626 );
nor ( w628 , w627 , g10 );
and ( w629 , w628 , g4 );
and ( w630 , g10 , w956 );
not ( w631 , w630 );
and ( w632 , w631 , g1 );
and ( w633 , w632 , w280 );
and ( w634 , w633 , g2 );
not ( w635 , w242 );
and ( w636 , w635 , w626 );
and ( w637 , w636 , w7213 );
nor ( w638 , w637 , g12 );
nor ( w639 , w638 , g3 );
and ( w640 , w639 , g11 );
nor ( w641 , w634 , w640 );
and ( w642 , w641 , w3 );
not ( w643 , w642 );
and ( w644 , w643 , w280 );
nor ( w645 , g1 , w89 );
and ( w646 , w12 , w3795 );
not ( w647 , w646 );
and ( w648 , w645 , w647 );
and ( w649 , w648 , w3 );
nor ( w650 , g1 , w231 );
nor ( w651 , w649 , w650 );
and ( w652 , w651 , g10 );
and ( w653 , w234 , g1 );
nor ( w654 , w653 , w83 );
nor ( w655 , w654 , w3 );
and ( w656 , w655 , g12 );
nor ( w657 , w44 , w656 );
nor ( w658 , w657 , g10 );
and ( w659 , w658 , g12 );
nor ( w660 , w652 , w659 );
nor ( w661 , w660 , w15 );
nor ( w662 , w661 , w264 );
nor ( w663 , w13 , w234 );
and ( w664 , w1898 , g1 );
nor ( w665 , w664 , w15 );
nor ( w666 , w649 , w47 );
and ( w667 , w666 , g13 );
and ( w668 , w667 , w5796 );
not ( w669 , w668 );
and ( w670 , w669 , w15 );
nor ( w671 , w665 , w670 );
not ( w672 , w671 );
and ( w673 , w672 , g10 );
and ( w674 , w6945 , w15 );
not ( w675 , w674 );
and ( w676 , w675 , w13 );
not ( w677 , w676 );
and ( w678 , w677 , w3 );
nor ( w679 , w674 , w527 );
not ( w680 , w679 );
and ( w681 , w680 , w8 );
nor ( w682 , w678 , w681 );
nor ( w683 , w682 , g4 );
and ( w684 , w6997 , w683 );
nor ( w685 , w673 , w684 );
nor ( w686 , w685 , g4 );
and ( w687 , w650 , w5796 );
not ( w688 , w687 );
and ( w689 , w688 , w15 );
nor ( w690 , w689 , w3 );
not ( w691 , w690 );
and ( w692 , w691 , g10 );
and ( w693 , w692 , w1025 );
nor ( w694 , w686 , w693 );
not ( w695 , w662 );
and ( w696 , w695 , w694 );
and ( w697 , w83 , w7183 );
nor ( w698 , w697 , w258 );
and ( w699 , w150 , g13 );
and ( w700 , w699 , w6997 );
and ( w701 , w700 , g4 );
nor ( w702 , w701 , w229 );
not ( w703 , w702 );
and ( w704 , w703 , g1 );
and ( w705 , w704 , g12 );
not ( w706 , w705 );
and ( w707 , w698 , w706 );
not ( w708 , w707 );
and ( w709 , w708 , g12 );
and ( w710 , w709 , w7097 );
nor ( w711 , w696 , w710 );
not ( w712 , w711 );
and ( w713 , w712 , g12 );
and ( w714 , w713 , w7097 );
not ( w715 , w714 );
and ( w716 , w715 , g11 );
and ( w717 , w6945 , w716 );
and ( w718 , w717 , g10 );
nor ( w719 , w718 , g2 );
and ( w720 , w719 , w626 );
and ( w721 , w720 , w6794 );
and ( w722 , w721 , w7183 );
and ( w723 , w47 , w15 );
and ( w724 , w723 , w7102 );
nor ( w725 , w724 , g12 );
not ( w726 , w725 );
and ( w727 , w726 , g11 );
and ( w728 , w727 , g2 );
and ( w729 , g1 , w473 );
not ( w730 , w729 );
and ( w731 , w730 , g10 );
not ( w732 , w731 );
and ( w733 , w732 , w626 );
nor ( w734 , w728 , w733 );
not ( w735 , w734 );
and ( w736 , w735 , g13 );
and ( w737 , w15 , w13 );
nor ( w738 , w737 , w9 );
not ( w739 , w738 );
and ( w740 , w739 , g2 );
nor ( w741 , w740 , w626 );
nor ( w742 , w741 , g10 );
and ( w743 , w742 , w6471 );
nor ( w744 , w743 , g12 );
nor ( w745 , w744 , g3 );
and ( w746 , w745 , g11 );
and ( w747 , w746 , w6945 );
and ( w748 , g2 , w3 );
and ( w749 , w4553 , g10 );
nor ( w750 , w748 , w626 );
nor ( w751 , w750 , g10 );
and ( w752 , w751 , w7102 );
and ( w753 , w752 , w7097 );
and ( w754 , w753 , g11 );
nor ( w755 , w749 , w754 );
nor ( w756 , w755 , w15 );
and ( w757 , w626 , w6997 );
not ( w758 , w757 );
and ( w759 , w758 , w3 );
nor ( w760 , w759 , w8 );
and ( w761 , w6997 , w603 );
not ( w762 , w761 );
and ( w763 , w762 , w8 );
nor ( w764 , w763 , w3 );
and ( w765 , w764 , w7102 );
nor ( w766 , w760 , w765 );
not ( w767 , w756 );
and ( w768 , w767 , w766 );
and ( w769 , w768 , w956 );
not ( w770 , w769 );
and ( w771 , w770 , g1 );
and ( w772 , w771 , w7102 );
and ( w773 , w772 , w7097 );
and ( w774 , w773 , g11 );
nor ( w775 , w747 , w774 );
nor ( w776 , w775 , g13 );
and ( w777 , w776 , w7102 );
nor ( w778 , w777 , g12 );
not ( w779 , w736 );
and ( w780 , w779 , w778 );
nor ( w781 , w780 , g3 );
and ( w782 , w781 , g11 );
nor ( w783 , w722 , w782 );
not ( w784 , w783 );
and ( w785 , w784 , g13 );
not ( w786 , w785 );
and ( w787 , w786 , w778 );
nor ( w788 , w787 , g4 );
nor ( w789 , w788 , g12 );
nor ( w790 , w789 , g3 );
and ( w791 , w790 , g11 );
nor ( w792 , w160 , w791 );
nor ( w793 , w792 , w3 );
and ( w794 , w793 , w7183 );
nor ( w795 , w794 , w782 );
not ( w796 , w795 );
and ( w797 , w796 , g13 );
not ( w798 , w797 );
and ( w799 , w798 , w778 );
nor ( w800 , w799 , g4 );
nor ( w801 , w800 , g12 );
nor ( w802 , w801 , g3 );
and ( w803 , w802 , g11 );
nor ( w804 , w644 , w803 );
nor ( w805 , w804 , w15 );
nor ( w806 , w805 , w782 );
not ( w807 , w806 );
and ( w808 , w807 , g13 );
not ( w809 , w808 );
and ( w810 , w809 , w778 );
nor ( w811 , w810 , g4 );
nor ( w812 , w811 , g12 );
nor ( w813 , w812 , g3 );
and ( w814 , w813 , g11 );
nor ( w815 , w629 , w814 );
and ( w816 , w815 , w6380 );
nor ( w817 , w816 , g3 );
and ( w818 , w817 , g11 );
and ( w819 , w525 , w818 );
and ( w820 , w819 , w6997 );
nor ( w821 , w86 , w820 );
not ( w822 , w821 );
and ( w823 , w822 , g4 );
and ( w824 , g12 , g13 );
and ( w825 , w824 , g1 );
not ( w826 , w825 );
and ( w827 , g1 , w826 );
and ( w828 , w827 , w7213 );
and ( w829 , w6380 , g2 );
not ( w830 , w829 );
and ( w831 , w830 , w13 );
and ( w832 , w831 , g11 );
and ( w833 , w832 , w7183 );
and ( w834 , w833 , w6997 );
not ( w835 , w828 );
and ( w836 , w835 , w834 );
and ( w837 , w836 , g3 );
and ( w838 , w473 , g11 );
and ( w839 , w838 , g1 );
and ( w840 , w543 , w7097 );
and ( w841 , w840 , g4 );
nor ( w842 , w839 , w841 );
not ( w843 , w842 );
and ( w844 , w843 , g4 );
not ( w845 , w234 );
and ( w846 , w845 , g13 );
nor ( w847 , w846 , w3 );
not ( w848 , w157 );
and ( w849 , w847 , w848 );
and ( w850 , w157 , w6997 );
nor ( w851 , w850 , g4 );
and ( w852 , w851 , w15 );
nor ( w853 , w849 , w852 );
nor ( w854 , w853 , w3 );
and ( w855 , w854 , g11 );
and ( w856 , w855 , w15 );
nor ( w857 , w62 , w856 );
not ( w858 , w857 );
and ( w859 , w858 , g11 );
and ( w860 , w859 , g2 );
and ( w861 , w95 , w7213 );
and ( w862 , w861 , w6997 );
and ( w863 , w862 , w13 );
nor ( w864 , g4 , w405 );
and ( w865 , w864 , w6471 );
nor ( w866 , w157 , g4 );
not ( w867 , w866 );
and ( w868 , w867 , g3 );
and ( w869 , w868 , w1025 );
and ( w870 , w869 , w6997 );
not ( w871 , w865 );
and ( w872 , w871 , w870 );
not ( w873 , w872 );
and ( w874 , w873 , g3 );
and ( w875 , w874 , w15 );
and ( w876 , w875 , w6794 );
and ( w877 , w876 , g11 );
nor ( w878 , w863 , w877 );
not ( w879 , w878 );
and ( w880 , w879 , g11 );
and ( w881 , w880 , w7213 );
and ( w882 , w881 , w6945 );
not ( w883 , w202 );
and ( w884 , w883 , g4 );
and ( w885 , w884 , g2 );
and ( w886 , w1 , g2 );
and ( w887 , w7097 , g4 );
nor ( w888 , w153 , g4 );
nor ( w889 , w887 , w888 );
nor ( w890 , w889 , g2 );
and ( w891 , w890 , w15 );
nor ( w892 , w886 , w891 );
nor ( w893 , w892 , g11 );
and ( w894 , w893 , g1 );
and ( w895 , w894 , w6794 );
and ( w896 , w895 , w15 );
and ( w897 , w896 , w6997 );
nor ( w898 , w44 , w897 );
nor ( w899 , w898 , g11 );
and ( w900 , w899 , w15 );
and ( w901 , w900 , w6997 );
and ( w902 , w901 , w7102 );
nor ( w903 , w902 , w897 );
and ( w904 , w903 , w1343 );
nor ( w905 , w904 , g2 );
and ( w906 , w905 , w15 );
and ( w907 , w906 , w6997 );
nor ( w908 , w885 , w907 );
not ( w909 , w908 );
and ( w910 , w909 , g1 );
and ( w911 , w910 , w3795 );
and ( w912 , w6161 , g2 );
not ( w913 , w912 );
and ( w914 , w913 , g4 );
nor ( w915 , w914 , w157 );
and ( w916 , w915 , g3 );
and ( w917 , w694 , w7102 );
and ( w918 , w917 , w7213 );
and ( w919 , w918 , w6794 );
and ( w920 , w919 , w15 );
nor ( w921 , w484 , w920 );
nor ( w922 , w921 , g3 );
and ( w923 , w922 , w6794 );
and ( w924 , w923 , w15 );
and ( w925 , w924 , w6997 );
nor ( w926 , w916 , w925 );
and ( w927 , w926 , w956 );
not ( w928 , w927 );
and ( w929 , w928 , g11 );
not ( w930 , w929 );
and ( w931 , w930 , g12 );
not ( w932 , w931 );
and ( w933 , w932 , g1 );
and ( w934 , w933 , w6794 );
and ( w935 , w934 , w15 );
and ( w936 , w935 , w6997 );
and ( w937 , g12 , w936 );
not ( w938 , w870 );
and ( w939 , w938 , g3 );
and ( w940 , w939 , w15 );
nor ( w941 , w937 , w940 );
not ( w942 , w850 );
and ( w943 , w942 , g3 );
nor ( w944 , g2 , w920 );
nor ( w945 , w944 , g3 );
and ( w946 , w945 , w6794 );
and ( w947 , w946 , w15 );
nor ( w948 , w943 , w947 );
nor ( w949 , w948 , g4 );
and ( w950 , w949 , g11 );
and ( w951 , w950 , g1 );
and ( w952 , w951 , w6794 );
and ( w953 , w952 , w15 );
not ( w954 , w953 );
and ( w955 , w941 , w954 );
not ( w956 , w473 );
and ( w957 , w955 , w956 );
not ( w958 , w957 );
and ( w959 , w958 , g11 );
nor ( w960 , w959 , w897 );
not ( w961 , w960 );
and ( w962 , w961 , g1 );
and ( w963 , w962 , w6794 );
and ( w964 , w963 , w15 );
and ( w965 , w964 , w6997 );
nor ( w966 , w911 , w965 );
not ( w967 , w966 );
and ( w968 , w967 , g3 );
and ( w969 , w901 , g2 );
nor ( w970 , w969 , w897 );
not ( w971 , w970 );
and ( w972 , w971 , g4 );
nor ( w973 , w44 , w965 );
nor ( w974 , w973 , g2 );
and ( w975 , w974 , w15 );
and ( w976 , w975 , w6997 );
nor ( w977 , w897 , w976 );
nor ( w978 , w977 , g4 );
and ( w979 , w978 , w7094 );
nor ( w980 , w972 , w979 );
and ( w981 , w531 , g4 );
nor ( w982 , g13 , g4 );
and ( w983 , w982 , g2 );
and ( w984 , w983 , w6997 );
nor ( w985 , w981 , w984 );
not ( w986 , w985 );
and ( w987 , w986 , g2 );
nor ( w988 , w554 , w555 );
nor ( w989 , w988 , g2 );
nor ( w990 , w989 , g12 );
not ( w991 , w987 );
and ( w992 , w991 , w990 );
and ( w993 , w992 , w3 );
not ( w994 , w993 );
and ( w995 , w994 , w280 );
and ( w996 , w540 , g2 );
and ( w997 , w574 , w7213 );
and ( w998 , w997 , w6794 );
and ( w999 , w998 , w15 );
nor ( w1000 , w996 , w999 );
not ( w1001 , w1000 );
and ( w1002 , w1001 , g4 );
and ( w1003 , w791 , w525 );
not ( w1004 , w145 );
and ( w1005 , g12 , w1004 );
not ( w1006 , w427 );
and ( w1007 , w1005 , w1006 );
nor ( w1008 , w1007 , g10 );
and ( w1009 , g12 , w1008 );
nor ( w1010 , w1009 , w965 );
not ( w1011 , w1003 );
and ( w1012 , w1011 , w1010 );
nor ( w1013 , w1012 , g10 );
nor ( w1014 , w1013 , g12 );
nor ( w1015 , w120 , g1 );
nor ( w1016 , w491 , w494 );
nor ( w1017 , w1016 , w473 );
not ( w1018 , w1017 );
and ( w1019 , w1018 , g1 );
nor ( w1020 , w1015 , w1019 );
and ( w1021 , w1020 , w3 );
nor ( w1022 , w965 , w145 );
not ( w1023 , w111 );
and ( w1024 , w1022 , w1023 );
not ( w1025 , w13 );
and ( w1026 , w1024 , w1025 );
and ( w1027 , w1026 , w1181 );
nor ( w1028 , w1027 , g10 );
not ( w1029 , w1021 );
and ( w1030 , w1029 , w1028 );
and ( w1031 , w1030 , g4 );
and ( w1032 , g2 , w6945 );
nor ( w1033 , w1032 , w1019 );
and ( w1034 , w1033 , w3 );
not ( w1035 , w1034 );
and ( w1036 , w1035 , w280 );
nor ( w1037 , w1008 , w965 );
and ( w1038 , w1037 , w1181 );
not ( w1039 , w1036 );
and ( w1040 , w1039 , w1038 );
nor ( w1041 , w1040 , g4 );
not ( w1042 , w1041 );
and ( w1043 , w1042 , g12 );
not ( w1044 , w1043 );
and ( w1045 , w1044 , g11 );
and ( w1046 , w1045 , w7097 );
and ( w1047 , w1046 , w15 );
and ( w1048 , w1047 , w6997 );
nor ( w1049 , w1031 , w1048 );
and ( w1050 , w1049 , g12 );
not ( w1051 , w1050 );
and ( w1052 , w1051 , g11 );
nor ( w1053 , w1052 , w820 );
nor ( w1054 , w1053 , g3 );
and ( w1055 , w1054 , w15 );
and ( w1056 , w1055 , w6997 );
not ( w1057 , w1014 );
and ( w1058 , w1057 , w1056 );
nor ( w1059 , w1058 , w820 );
not ( w1060 , w1002 );
and ( w1061 , w1060 , w1059 );
nor ( w1062 , w1061 , w3 );
and ( w1063 , w1062 , w1056 );
nor ( w1064 , w1063 , w820 );
not ( w1065 , w1064 );
and ( w1066 , w1065 , w15 );
nor ( w1067 , w995 , w1066 );
and ( w1068 , w1067 , w6380 );
not ( w1069 , w1068 );
and ( w1070 , w1069 , w1056 );
not ( w1071 , w1070 );
and ( w1072 , w980 , w1071 );
and ( w1073 , w1072 , w1181 );
nor ( w1074 , w1073 , g3 );
and ( w1075 , w1074 , w15 );
nor ( w1076 , w968 , w1075 );
not ( w1077 , w1076 );
and ( w1078 , w1077 , w15 );
and ( w1079 , w1078 , w6997 );
nor ( w1080 , w882 , w1079 );
not ( w1081 , w1080 );
and ( w1082 , w1081 , g3 );
nor ( w1083 , w1082 , w1075 );
not ( w1084 , w1083 );
and ( w1085 , w1084 , w15 );
and ( w1086 , w1085 , w6997 );
nor ( w1087 , w860 , w1086 );
nor ( w1088 , w1087 , g1 );
nor ( w1089 , w1088 , w1079 );
not ( w1090 , w1089 );
and ( w1091 , w1090 , g3 );
nor ( w1092 , w1091 , w1075 );
not ( w1093 , w1092 );
and ( w1094 , w1093 , w15 );
and ( w1095 , w1094 , w6997 );
nor ( w1096 , w839 , w1095 );
not ( w1097 , w844 );
and ( w1098 , w1097 , w1096 );
not ( w1099 , w1098 );
and ( w1100 , w1099 , g2 );
nor ( w1101 , w220 , g13 );
and ( w1102 , w1101 , g4 );
not ( w1103 , w1102 );
and ( w1104 , w1103 , w1096 );
not ( w1105 , w1104 );
and ( w1106 , w1105 , g3 );
and ( w1107 , w1106 , w7213 );
nor ( w1108 , w82 , w659 );
nor ( w1109 , w1108 , g3 );
and ( w1110 , w1109 , g11 );
not ( w1111 , w1110 );
and ( w1112 , g12 , w1111 );
not ( w1113 , w1112 );
and ( w1114 , w1113 , g1 );
nor ( w1115 , w1114 , w1095 );
not ( w1116 , w1115 );
and ( w1117 , w1116 , g4 );
nor ( w1118 , w1117 , w820 );
nor ( w1119 , w1118 , g3 );
and ( w1120 , w1119 , w7213 );
not ( w1121 , w1120 );
and ( w1122 , w1121 , w8 );
nor ( w1123 , w1122 , w3 );
and ( w1124 , w1123 , g11 );
and ( w1125 , w1124 , w7183 );
nor ( w1126 , w1125 , w1095 );
nor ( w1127 , w1126 , g10 );
nor ( w1128 , w1107 , w1127 );
and ( w1129 , w1128 , w8 );
nor ( w1130 , w1129 , w3 );
and ( w1131 , w1130 , g11 );
and ( w1132 , w1131 , w7183 );
nor ( w1133 , w1132 , w1095 );
nor ( w1134 , w1133 , g10 );
nor ( w1135 , w1100 , w1134 );
and ( w1136 , w1135 , w8 );
nor ( w1137 , w1136 , w3 );
and ( w1138 , w1137 , g11 );
and ( w1139 , w1138 , w7183 );
nor ( w1140 , w1139 , w1095 );
nor ( w1141 , w1140 , g10 );
nor ( w1142 , w634 , w839 );
nor ( w1143 , w1142 , g3 );
and ( w1144 , w1143 , w7102 );
and ( w1145 , w1144 , g11 );
nor ( w1146 , w1141 , w1145 );
and ( w1147 , w1146 , w1181 );
nor ( w1148 , w1147 , g3 );
and ( w1149 , w1148 , w7102 );
and ( w1150 , w1149 , w280 );
nor ( w1151 , w1150 , w1141 );
nor ( w1152 , w1151 , w15 );
nor ( w1153 , w1152 , w1095 );
not ( w1154 , w837 );
and ( w1155 , w1154 , w1153 );
nor ( w1156 , w1155 , g4 );
and ( w1157 , w1156 , w280 );
nor ( w1158 , w1157 , w1141 );
not ( w1159 , w823 );
and ( w1160 , w1159 , w1158 );
not ( w1161 , w1160 );
and ( w1162 , w1161 , w280 );
nor ( w1163 , w1162 , w1141 );
not ( w1164 , w1163 );
and ( w1165 , w1164 , g11 );
and ( w1166 , w1165 , w7183 );
nor ( w1167 , w1166 , w1095 );
nor ( w1168 , w1167 , g10 );
nor ( w1169 , w1168 , g2 );
and ( w1170 , w1169 , w6380 );
not ( w1171 , w531 );
and ( w1172 , w1171 , g2 );
nor ( w1173 , w1172 , g3 );
and ( w1174 , w1173 , g1 );
and ( w1175 , w1174 , g4 );
and ( w1176 , w1175 , w7183 );
nor ( w1177 , w1176 , w1095 );
nor ( w1178 , w1177 , g10 );
nor ( w1179 , w370 , w1178 );
and ( w1180 , w1179 , w6380 );
not ( w1181 , w820 );
and ( w1182 , w1181 , g2 );
and ( w1183 , w1182 , g12 );
nor ( w1184 , w1183 , w15 );
nor ( w1185 , w1184 , w1095 );
nor ( w1186 , w1185 , g10 );
not ( w1187 , w1180 );
and ( w1188 , w1187 , w1186 );
and ( w1189 , w1188 , g1 );
nor ( w1190 , w1189 , w839 );
not ( w1191 , w1190 );
and ( w1192 , w1191 , g4 );
and ( w1193 , w1192 , g11 );
and ( w1194 , w1193 , w7183 );
nor ( w1195 , w1194 , w1095 );
nor ( w1196 , w1195 , g10 );
not ( w1197 , w1196 );
and ( w1198 , w1169 , w1197 );
not ( w1199 , w1198 );
and ( w1200 , w1199 , g4 );
not ( w1201 , w1200 );
and ( w1202 , w1201 , w1158 );
not ( w1203 , w1202 );
and ( w1204 , w1203 , w280 );
nor ( w1205 , w1204 , w1141 );
nor ( w1206 , w1205 , w15 );
nor ( w1207 , w1206 , w1095 );
nor ( w1208 , w1207 , g10 );
not ( w1209 , w1208 );
and ( w1210 , w1209 , g12 );
nor ( w1211 , w1210 , g1 );
nor ( w1212 , w1211 , w1196 );
not ( w1213 , w1212 );
and ( w1214 , w1213 , g4 );
not ( w1215 , w1214 );
and ( w1216 , w1215 , w1158 );
not ( w1217 , w1216 );
and ( w1218 , w1217 , w280 );
nor ( w1219 , w1218 , w1141 );
not ( w1220 , w1219 );
and ( w1221 , w1220 , g11 );
and ( w1222 , w1221 , w7183 );
nor ( w1223 , w1222 , w1095 );
nor ( w1224 , w1223 , g10 );
not ( w1225 , w1170 );
and ( w1226 , w1225 , w1224 );
nor ( w1227 , w1226 , w1196 );
not ( w1228 , w77 );
and ( w1229 , w1228 , w1227 );
and ( w1230 , w6997 , w1229 );
nor ( w1231 , w1230 , g11 );
nor ( w1232 , w1231 , w839 );
and ( w1233 , w1281 , g1 );
not ( w1234 , w1233 );
and ( w1235 , w1229 , w1234 );
nor ( w1236 , w1235 , w3 );
nor ( w1237 , w1236 , w13 );
nor ( w1238 , w1237 , w1230 );
and ( w1239 , w1238 , g4 );
and ( w1240 , w6945 , w1229 );
nor ( w1241 , w1240 , w1230 );
and ( w1242 , w1241 , w6794 );
not ( w1243 , w1242 );
and ( w1244 , w1243 , w1229 );
nor ( w1245 , g13 , w1230 );
not ( w1246 , w1245 );
and ( w1247 , w1246 , w1229 );
not ( w1248 , w1247 );
and ( w1249 , w1248 , w13 );
not ( w1250 , w1249 );
and ( w1251 , w1250 , w1229 );
and ( w1252 , w1251 , w1343 );
not ( w1253 , w1252 );
and ( w1254 , w1253 , g11 );
not ( w1255 , w1254 );
and ( w1256 , w1244 , w1255 );
nor ( w1257 , w1256 , g4 );
not ( w1258 , w1257 );
and ( w1259 , w1258 , w1229 );
nor ( w1260 , w1259 , w15 );
not ( w1261 , w1260 );
and ( w1262 , w1261 , w1229 );
and ( w1263 , w1262 , w7097 );
nor ( w1264 , w1263 , w1230 );
nor ( w1265 , w1239 , w1264 );
nor ( w1266 , w1265 , w15 );
and ( w1267 , g11 , w1343 );
and ( w1268 , w1267 , w1229 );
nor ( w1269 , w1268 , w1230 );
not ( w1270 , w1269 );
and ( w1271 , w1270 , w3 );
and ( w1272 , w1229 , w7183 );
and ( w1273 , w1272 , g4 );
and ( w1274 , w1229 , w7102 );
nor ( w1275 , w1273 , w1274 );
nor ( w1276 , w292 , w1230 );
not ( w1277 , w1276 );
and ( w1278 , w1277 , g4 );
nor ( w1279 , w1278 , w1230 );
and ( w1280 , w1279 , w7183 );
not ( w1281 , w1232 );
and ( w1282 , w1281 , w15 );
nor ( w1283 , w1282 , g2 );
nor ( w1284 , w1283 , w1230 );
nor ( w1285 , w1284 , g3 );
nor ( w1286 , w1285 , w1230 );
nor ( w1287 , w1280 , w1286 );
and ( w1288 , w1287 , w1229 );
not ( w1289 , w1288 );
and ( w1290 , w1289 , g1 );
not ( w1291 , w1290 );
and ( w1292 , w1291 , w1229 );
and ( w1293 , w1292 , w3 );
not ( w1294 , w1293 );
and ( w1295 , w1294 , w280 );
nor ( w1296 , w1295 , g2 );
nor ( w1297 , w1296 , w1230 );
nor ( w1298 , w1297 , g3 );
nor ( w1299 , w1298 , w1230 );
nor ( w1300 , w1275 , w1299 );
nor ( w1301 , w1300 , w1230 );
not ( w1302 , w1301 );
and ( w1303 , w1302 , w3 );
not ( w1304 , w1303 );
and ( w1305 , w1304 , w13 );
nor ( w1306 , w686 , w1230 );
and ( w1307 , w234 , g10 );
not ( w1308 , w1306 );
and ( w1309 , w1308 , w1307 );
nor ( w1310 , w1309 , w1230 );
nor ( w1311 , w1310 , g2 );
nor ( w1312 , w1311 , w1230 );
nor ( w1313 , w1312 , g3 );
nor ( w1314 , w1313 , w1230 );
and ( w1315 , w1314 , g1 );
not ( w1316 , w1315 );
and ( w1317 , w1229 , w1316 );
and ( w1318 , w1317 , w7102 );
nor ( w1319 , w1318 , w1230 );
nor ( w1320 , w15 , w1319 );
nor ( w1321 , w1320 , w1230 );
and ( w1322 , w251 , w1391 );
nor ( w1323 , w1322 , w236 );
and ( w1324 , w1323 , w1229 );
not ( w1325 , w1324 );
and ( w1326 , w1325 , w15 );
not ( w1327 , w1326 );
and ( w1328 , w1327 , w1229 );
nor ( w1329 , w1328 , w3 );
not ( w1330 , w1329 );
and ( w1331 , w1330 , w1229 );
and ( w1332 , w1331 , w7213 );
nor ( w1333 , w1332 , w1230 );
nor ( w1334 , w1333 , g3 );
nor ( w1335 , w1334 , w1230 );
and ( w1336 , w1335 , g4 );
and ( w1337 , w1245 , w7102 );
nor ( w1338 , w1336 , w1337 );
nor ( w1339 , w1338 , g1 );
and ( w1340 , w1391 , g4 );
not ( w1341 , w1340 );
and ( w1342 , w1341 , w1229 );
not ( w1343 , w839 );
and ( w1344 , w1342 , w1343 );
not ( w1345 , w1344 );
and ( w1346 , w1345 , g1 );
and ( w1347 , w1346 , g11 );
nor ( w1348 , w1347 , g3 );
not ( w1349 , w1339 );
and ( w1350 , w1349 , w1348 );
not ( w1351 , w1350 );
and ( w1352 , w1351 , g11 );
and ( w1353 , w1352 , w1391 );
and ( w1354 , w1353 , w15 );
and ( w1355 , w1354 , w6794 );
nor ( w1356 , w1355 , g2 );
nor ( w1357 , w1356 , w1230 );
nor ( w1358 , w1357 , g3 );
and ( w1359 , w1229 , w1358 );
nor ( w1360 , w1359 , w1230 );
not ( w1361 , w1360 );
and ( w1362 , w15 , w1361 );
nor ( w1363 , w1362 , w1230 );
and ( w1364 , w1363 , w6794 );
not ( w1365 , w1364 );
and ( w1366 , w1365 , w1229 );
and ( w1367 , w1366 , w7213 );
nor ( w1368 , w1367 , w1230 );
nor ( w1369 , w1272 , w1230 );
and ( w1370 , w1401 , g2 );
and ( w1371 , w1229 , w15 );
and ( w1372 , w1371 , w7213 );
nor ( w1373 , w1370 , w1372 );
and ( w1374 , w1373 , w1391 );
not ( w1375 , w1374 );
and ( w1376 , w1375 , w3 );
nor ( w1377 , w9 , g2 );
and ( w1378 , w1377 , w1229 );
and ( w1379 , w1378 , w7183 );
nor ( w1380 , w1379 , w1230 );
nor ( w1381 , w1380 , w13 );
nor ( w1382 , w1376 , w1381 );
not ( w1383 , w1382 );
and ( w1384 , w1383 , g4 );
and ( w1385 , w1229 , g2 );
and ( w1386 , w1385 , w15 );
nor ( w1387 , w1386 , w1230 );
and ( w1388 , w1386 , w3 );
nor ( w1389 , w1388 , w1230 );
and ( w1390 , w1389 , w7094 );
not ( w1391 , w1230 );
and ( w1392 , g13 , w1391 );
and ( w1393 , w1392 , w6380 );
not ( w1394 , w1393 );
and ( w1395 , w1394 , g2 );
and ( w1396 , w1395 , w1229 );
and ( w1397 , w15 , w1396 );
nor ( w1398 , w1397 , w1230 );
not ( w1399 , w1398 );
and ( w1400 , w1399 , w3 );
not ( w1401 , w1369 );
and ( w1402 , w1401 , g4 );
nor ( w1403 , w15 , w1230 );
not ( w1404 , w1403 );
and ( w1405 , w1404 , w1229 );
and ( w1406 , w1405 , w7102 );
nor ( w1407 , w1402 , w1406 );
nor ( w1408 , w1407 , w13 );
nor ( w1409 , w1400 , w1408 );
nor ( w1410 , w1409 , w839 );
not ( w1411 , w1410 );
and ( w1412 , w1411 , g11 );
and ( w1413 , w1412 , g1 );
nor ( w1414 , w1390 , w1413 );
not ( w1415 , w1414 );
and ( w1416 , w1415 , g1 );
not ( w1417 , w1416 );
and ( w1418 , w1417 , w1229 );
not ( w1419 , w1387 );
and ( w1420 , w1419 , w1418 );
and ( w1421 , w1420 , w7102 );
nor ( w1422 , w1384 , w1421 );
and ( w1423 , w1368 , w1422 );
nor ( w1424 , w1423 , g3 );
nor ( w1425 , w1424 , w1230 );
and ( w1426 , w1321 , w1425 );
and ( w1427 , w1426 , w6794 );
not ( w1428 , w1427 );
and ( w1429 , w1428 , w1229 );
and ( w1430 , w1429 , w7213 );
nor ( w1431 , w1430 , w1230 );
and ( w1432 , w1431 , w1422 );
nor ( w1433 , w1432 , g3 );
nor ( w1434 , w1433 , w1230 );
nor ( w1435 , w1305 , w1434 );
and ( w1436 , w1435 , w7213 );
not ( w1437 , w1436 );
and ( w1438 , w1437 , w1422 );
nor ( w1439 , w1438 , g3 );
nor ( w1440 , w1230 , w1439 );
not ( w1441 , w1271 );
and ( w1442 , w1441 , w1440 );
and ( w1443 , w1442 , g1 );
not ( w1444 , w1443 );
and ( w1445 , w1444 , g4 );
and ( w1446 , w1445 , g2 );
nor ( w1447 , w1446 , w1439 );
nor ( w1448 , w1447 , g3 );
and ( w1449 , w1229 , w1448 );
nor ( w1450 , w1449 , w1230 );
not ( w1451 , w1450 );
and ( w1452 , w1451 , g4 );
nor ( w1453 , w1452 , w1230 );
and ( w1454 , w1453 , w15 );
not ( w1455 , w1454 );
and ( w1456 , w1455 , w1229 );
and ( w1457 , w1456 , g2 );
nor ( w1458 , w1457 , w1230 );
and ( w1459 , w1458 , w1466 );
and ( w1460 , w1459 , w1422 );
nor ( w1461 , w1460 , g3 );
nor ( w1462 , w1461 , w1230 );
nor ( w1463 , w1266 , w1462 );
and ( w1464 , w1463 , g2 );
nor ( w1465 , w1464 , w1230 );
not ( w1466 , w1439 );
and ( w1467 , w1465 , w1466 );
and ( w1468 , w1467 , w6945 );
and ( w1469 , w1233 , w1467 );
and ( w1470 , w1469 , g2 );
and ( w1471 , w1470 , g4 );
and ( w1472 , w1469 , w7213 );
and ( w1473 , w1472 , w7102 );
and ( w1474 , w7097 , w1467 );
nor ( w1475 , w1473 , w1474 );
and ( w1476 , w1475 , w1229 );
nor ( w1477 , w1476 , w15 );
and ( w1478 , w1467 , g2 );
and ( w1479 , w1478 , w7102 );
nor ( w1480 , w1479 , w1474 );
and ( w1481 , w1480 , w1229 );
not ( w1482 , w1481 );
and ( w1483 , w1482 , w15 );
nor ( w1484 , w1477 , w1483 );
not ( w1485 , w1484 );
and ( w1486 , w1485 , w13 );
and ( w1487 , w1467 , w7213 );
nor ( w1488 , w1487 , w1474 );
and ( w1489 , w1488 , w1229 );
nor ( w1490 , w1489 , w15 );
nor ( w1491 , w1490 , w1474 );
and ( w1492 , w1491 , w1229 );
not ( w1493 , w1492 );
and ( w1494 , w1493 , g4 );
nor ( w1495 , w1494 , w1474 );
nor ( w1496 , w1495 , w3 );
nor ( w1497 , w1470 , w1474 );
and ( w1498 , w1497 , w1229 );
nor ( w1499 , w1498 , w15 );
not ( w1500 , w1474 );
and ( w1501 , w1500 , w1229 );
not ( w1502 , w1499 );
and ( w1503 , w1502 , w1501 );
and ( w1504 , w1472 , w15 );
not ( w1505 , w1504 );
and ( w1506 , w1503 , w1505 );
nor ( w1507 , w1506 , g4 );
and ( w1508 , w1507 , w6794 );
not ( w1509 , w1508 );
and ( w1510 , w1509 , w1501 );
not ( w1511 , w1496 );
and ( w1512 , w1511 , w1510 );
nor ( w1513 , w1512 , g11 );
nor ( w1514 , w1513 , w839 );
not ( w1515 , w1514 );
and ( w1516 , w1515 , g1 );
not ( w1517 , w1516 );
and ( w1518 , w1517 , w1501 );
not ( w1519 , w1486 );
and ( w1520 , w1519 , w1518 );
nor ( w1521 , w1520 , g11 );
nor ( w1522 , w1521 , w839 );
not ( w1523 , w1522 );
and ( w1524 , w1523 , g1 );
not ( w1525 , w1524 );
and ( w1526 , w1525 , w1501 );
not ( w1527 , w1471 );
and ( w1528 , w1527 , w1526 );
not ( w1529 , w1528 );
and ( w1530 , w1529 , w1467 );
and ( w1531 , w1530 , w7183 );
nor ( w1532 , w1531 , w1483 );
not ( w1533 , w1532 );
and ( w1534 , w1533 , w13 );
not ( w1535 , w1534 );
and ( w1536 , w1535 , w1518 );
nor ( w1537 , w1536 , g11 );
nor ( w1538 , w1537 , w839 );
not ( w1539 , w1538 );
and ( w1540 , w1539 , g1 );
not ( w1541 , w1540 );
and ( w1542 , w1541 , w1501 );
not ( w1543 , w1468 );
and ( w1544 , w1543 , w1542 );
not ( w1545 , w1544 );
and ( w1546 , w1545 , w1467 );
not ( w1547 , w1546 );
and ( w1548 , w1547 , w3 );
not ( w1549 , w1548 );
and ( w1550 , w1549 , w280 );
nor ( w1551 , w1550 , w1474 );
nor ( w1552 , w1551 , w15 );
and ( w1553 , w1467 , g1 );
not ( w1554 , w1553 );
and ( w1555 , w1554 , w1542 );
not ( w1556 , w1555 );
and ( w1557 , w1556 , w1467 );
and ( w1558 , w1557 , w15 );
nor ( w1559 , w1558 , w1474 );
and ( w1560 , w1559 , w1501 );
not ( w1561 , w1552 );
and ( w1562 , w1561 , w1560 );
and ( w1563 , w1562 , w1542 );
not ( w1564 , w1563 );
and ( w1565 , w1564 , g4 );
not ( w1566 , w1565 );
and ( w1567 , w1566 , w1542 );
and ( w1568 , w1468 , g11 );
not ( w1569 , w1568 );
and ( w1570 , w1569 , w1542 );
not ( w1571 , w1570 );
and ( w1572 , w1571 , w1467 );
and ( w1573 , w1572 , w6794 );
not ( w1574 , w1573 );
and ( w1575 , w1574 , w1229 );
and ( w1576 , w1575 , w1501 );
and ( w1577 , w1576 , w1542 );
nor ( w1578 , w1577 , w15 );
not ( w1579 , w1572 );
and ( w1580 , w1579 , w3 );
and ( w1581 , w1580 , w1542 );
not ( w1582 , w1581 );
and ( w1583 , w1582 , w1467 );
and ( w1584 , w1583 , w280 );
not ( w1585 , w1584 );
and ( w1586 , w1585 , w1542 );
not ( w1587 , w1586 );
and ( w1588 , w1587 , w15 );
and ( w1589 , w1588 , w1467 );
nor ( w1590 , w1589 , w1474 );
not ( w1591 , w1578 );
and ( w1592 , w1591 , w1590 );
not ( w1593 , w1592 );
and ( w1594 , w1593 , w1467 );
and ( w1595 , w1594 , w7102 );
not ( w1596 , w1595 );
and ( w1597 , w1596 , w1229 );
and ( w1598 , w1597 , w1501 );
and ( w1599 , w1598 , w1542 );
nor ( w1600 , w1599 , g2 );
nor ( w1601 , w1600 , w1474 );
and ( w1602 , w1567 , w1601 );
not ( w1603 , w1602 );
and ( w1604 , w1603 , w1467 );
and ( w1605 , w1604 , w7213 );
nor ( w1606 , w1605 , w1474 );
and ( w1607 , w7213 , w1606 );
nor ( w1608 , w1607 , w1230 );
and ( w1609 , w1468 , g13 );
and ( w1610 , w1606 , w1229 );
and ( w1611 , w1467 , w1608 );
and ( w1612 , w1611 , g1 );
nor ( w1613 , w1612 , w1474 );
and ( w1614 , w1613 , w1229 );
nor ( w1615 , w1614 , g4 );
not ( w1616 , w1615 );
and ( w1617 , w1616 , w1606 );
not ( w1618 , w1617 );
and ( w1619 , w1618 , w15 );
not ( w1620 , w1619 );
and ( w1621 , w1610 , w1620 );
nor ( w1622 , w1621 , w3 );
not ( w1623 , w1622 );
and ( w1624 , w1623 , w1542 );
and ( w1625 , w1624 , w1606 );
and ( w1626 , w1553 , g13 );
and ( w1627 , w1626 , w1611 );
not ( w1628 , w1627 );
and ( w1629 , w1628 , w1606 );
not ( w1630 , w1629 );
and ( w1631 , w1630 , g4 );
not ( w1632 , w1631 );
and ( w1633 , w1632 , w1606 );
not ( w1634 , w1633 );
and ( w1635 , w1634 , w15 );
nor ( w1636 , w1635 , w1474 );
and ( w1637 , w1636 , w1501 );
and ( w1638 , w1637 , w1542 );
not ( w1639 , w1638 );
and ( w1640 , w1639 , w1467 );
not ( w1641 , w1640 );
and ( w1642 , w1641 , w3 );
and ( w1643 , w1642 , w1542 );
not ( w1644 , w1643 );
and ( w1645 , w1644 , w13 );
not ( w1646 , w1645 );
and ( w1647 , w1646 , w1229 );
and ( w1648 , w1610 , w1542 );
and ( w1649 , w1647 , w1648 );
and ( w1650 , w1625 , w1649 );
not ( w1651 , w1609 );
and ( w1652 , w1651 , w1650 );
not ( w1653 , w1652 );
and ( w1654 , w1653 , w1611 );
not ( w1655 , w1654 );
and ( w1656 , w1655 , w3 );
not ( w1657 , w1656 );
and ( w1658 , w1657 , w1611 );
and ( w1659 , w1658 , w13 );
not ( w1660 , w1659 );
and ( w1661 , w1660 , w1229 );
and ( w1662 , w1661 , w1606 );
not ( w1663 , w1662 );
and ( w1664 , w1663 , g4 );
not ( w1665 , w1664 );
and ( w1666 , w1665 , w1606 );
and ( w1667 , w1666 , w1542 );
and ( w1668 , w1611 , w6945 );
not ( w1669 , w1668 );
and ( w1670 , w1669 , w1650 );
not ( w1671 , w1670 );
and ( w1672 , w1671 , w1611 );
and ( w1673 , w1672 , w6794 );
not ( w1674 , w1673 );
and ( w1675 , w1674 , w1606 );
and ( w1676 , w1675 , w1229 );
and ( w1677 , w1676 , w1648 );
nor ( w1678 , w1677 , g4 );
and ( w1679 , w1678 , w15 );
not ( w1680 , w1679 );
and ( w1681 , w1667 , w1680 );
not ( w1682 , w1681 );
and ( w1683 , w1682 , w1467 );
not ( w1684 , w1683 );
and ( w1685 , w15 , w1684 );
nor ( w1686 , w1685 , w1230 );
and ( w1687 , w1608 , w1686 );
and ( w1688 , w1687 , w1467 );
and ( w1689 , w1688 , g1 );
not ( w1690 , w1689 );
and ( w1691 , w1690 , w1650 );
not ( w1692 , w1691 );
and ( w1693 , w1692 , w1467 );
and ( w1694 , w1683 , w15 );
nor ( w1695 , w1694 , w1474 );
and ( w1696 , w1695 , w1501 );
not ( w1697 , w1693 );
and ( w1698 , w1697 , w1696 );
not ( w1699 , w1698 );
and ( w1700 , w1699 , w280 );
not ( w1701 , w1694 );
and ( w1702 , w1701 , w1606 );
and ( w1703 , w1702 , w1229 );
not ( w1704 , w1700 );
and ( w1705 , w1704 , w1703 );
and ( w1706 , w1705 , w1542 );
and ( w1707 , g1 , w1706 );
not ( w1708 , w1706 );
and ( w1709 , w1708 , w1467 );
and ( w1710 , w1709 , w7102 );
not ( w1711 , w1710 );
and ( w1712 , w1711 , w1606 );
and ( w1713 , w7102 , w1712 );
not ( w1714 , w1713 );
and ( w1715 , w1714 , w1467 );
and ( w1716 , w3 , w1706 );
not ( w1717 , w1716 );
and ( w1718 , w1715 , w1717 );
and ( w1719 , w1718 , w1688 );
not ( w1720 , w1707 );
and ( t_0 , w1720 , w1719 );
nor ( w1721 , g1 , g10 );
and ( w1722 , w231 , w7102 );
and ( w1723 , w1722 , g3 );
and ( w1724 , w982 , w7097 );
and ( w1725 , w1724 , w7183 );
and ( w1726 , w6794 , g7 );
nor ( w1727 , w1726 , w2 );
nor ( w1728 , w3 , w1727 );
nor ( w1729 , w12 , w1728 );
and ( w1730 , w12 , w3 );
nor ( w1731 , w228 , w1730 );
not ( w1732 , g5 );
and ( w1733 , g7 , w1732 );
nor ( w1734 , w12 , w1733 );
nor ( w1735 , g5 , w1733 );
nor ( w1736 , w1734 , w1735 );
nor ( w1737 , w1736 , w1730 );
nor ( w1738 , w1731 , w1737 );
not ( w1739 , w1738 );
and ( w1740 , w1728 , w1739 );
nor ( w1741 , w1740 , w15 );
nor ( w1742 , w1741 , w740 );
not ( w1743 , w1742 );
and ( w1744 , w1743 , g2 );
and ( w1745 , w1744 , g13 );
nor ( w1746 , g4 , g2 );
and ( w1747 , w1746 , w2357 );
and ( w1748 , w1747 , g13 );
and ( w1749 , w1748 , w15 );
and ( w1750 , w1749 , g12 );
and ( w1751 , w1750 , g11 );
and ( w1752 , w1751 , w7097 );
nor ( w1753 , w1745 , w1752 );
not ( w1754 , w1753 );
and ( w1755 , w1754 , g12 );
and ( w1756 , w1755 , g11 );
and ( w1757 , w1756 , w7097 );
and ( w1758 , w1757 , w7102 );
and ( w1759 , w231 , w7213 );
and ( w1760 , w1759 , w7102 );
and ( w1761 , w1760 , w7183 );
and ( w1762 , w1761 , g12 );
nor ( w1763 , w1762 , w1727 );
nor ( w1764 , w1763 , w1731 );
and ( w1765 , w1764 , g11 );
nor ( w1766 , w1758 , w1765 );
nor ( w1767 , w1766 , w15 );
and ( w1768 , w1767 , w2357 );
and ( w1769 , w1768 , w6997 );
and ( w1770 , w1758 , w6997 );
nor ( w1771 , w1769 , w1770 );
nor ( w1772 , w1771 , w15 );
and ( w1773 , w1772 , g2 );
nor ( w1774 , w477 , w1772 );
not ( w1775 , w1774 );
and ( w1776 , w1775 , g2 );
and ( w1777 , w1776 , w6471 );
and ( w1778 , w370 , w2606 );
and ( w1779 , w1778 , w2404 );
nor ( w1780 , w1751 , w1770 );
not ( w1781 , w1780 );
and ( w1782 , w1781 , w15 );
and ( w1783 , w1782 , w6997 );
nor ( w1784 , w1779 , w1783 );
not ( w1785 , w1770 );
and ( w1786 , w1784 , w1785 );
not ( w1787 , w1786 );
and ( w1788 , w1787 , g13 );
and ( w1789 , w1788 , w7102 );
and ( w1790 , w1789 , w15 );
and ( w1791 , w1790 , w6997 );
and ( w1792 , w1791 , g12 );
and ( w1793 , w1792 , g11 );
not ( w1794 , w1793 );
and ( w1795 , w1794 , w1737 );
and ( w1796 , g13 , g4 );
nor ( w1797 , w1796 , w1768 );
nor ( w1798 , w1797 , w15 );
and ( w1799 , w6471 , g3 );
not ( w1800 , w95 );
and ( w1801 , w1800 , g2 );
not ( w1802 , w1801 );
and ( w1803 , w1802 , g2 );
nor ( w1804 , w1746 , w1757 );
nor ( w1805 , w1804 , g4 );
not ( w1806 , w1805 );
and ( w1807 , w1806 , g12 );
not ( w1808 , w1807 );
and ( w1809 , w1808 , g11 );
nor ( w1810 , w92 , w1809 );
and ( w1811 , w699 , g12 );
and ( w1812 , w1811 , w6997 );
and ( w1813 , w1812 , g11 );
and ( w1814 , w1813 , w7213 );
nor ( w1815 , w1814 , g2 );
not ( w1816 , w1815 );
and ( w1817 , w1816 , g13 );
and ( w1818 , w1817 , g1 );
and ( w1819 , w1818 , g4 );
and ( w1820 , w1819 , w15 );
and ( w1821 , w1820 , w2357 );
and ( w1822 , w1821 , g12 );
and ( w1823 , w1822 , g11 );
nor ( w1824 , w1758 , w1823 );
and ( w1825 , w1824 , w2111 );
nor ( w1826 , w1825 , w1731 );
not ( w1827 , w1826 );
and ( w1828 , w1810 , w1827 );
and ( w1829 , w1828 , g13 );
and ( w1830 , w150 , g12 );
and ( w1831 , w1830 , w6997 );
and ( w1832 , w1831 , g11 );
not ( w1833 , w1832 );
and ( w1834 , w1833 , g3 );
not ( w1835 , w1834 );
and ( w1836 , w1835 , w15 );
and ( w1837 , w1836 , g11 );
and ( w1838 , w1837 , w7213 );
and ( w1839 , w1838 , w6471 );
and ( w1840 , w1839 , g4 );
and ( w1841 , w1840 , g12 );
and ( w1842 , w1841 , w2357 );
nor ( w1843 , w1842 , w1823 );
nor ( w1844 , w1843 , g2 );
nor ( w1845 , w1032 , w1844 );
and ( w1846 , w1845 , w6471 );
not ( w1847 , w1846 );
and ( w1848 , w1847 , w15 );
not ( w1849 , w1737 );
and ( w1850 , w1848 , w1849 );
and ( w1851 , w1850 , g11 );
not ( w1852 , w1829 );
and ( w1853 , w1852 , w1851 );
not ( w1854 , w1853 );
and ( w1855 , w1854 , g12 );
not ( w1856 , w1855 );
and ( w1857 , w1856 , w15 );
and ( w1858 , w1857 , w7097 );
nor ( w1859 , w1858 , g3 );
nor ( w1860 , w1859 , w1731 );
not ( w1861 , w1803 );
and ( w1862 , w1861 , w1860 );
not ( w1863 , w1862 );
and ( w1864 , w1863 , g12 );
not ( w1865 , w1864 );
and ( w1866 , w15 , w1865 );
nor ( w1867 , w1866 , g3 );
nor ( w1868 , w1867 , w1731 );
and ( w1869 , w1868 , g11 );
not ( w1870 , w1799 );
and ( w1871 , w1870 , w1869 );
and ( w1872 , w1871 , g2 );
and ( w1873 , w1837 , w1860 );
and ( w1874 , w1873 , w7213 );
and ( w1875 , w1874 , g4 );
and ( w1876 , w1875 , g12 );
nor ( w1877 , w1872 , w1876 );
and ( w1878 , w1826 , w15 );
not ( w1879 , w1878 );
and ( w1880 , w1877 , w1879 );
not ( w1881 , w1880 );
and ( w1882 , w1881 , g4 );
nor ( w1883 , w1882 , w1751 );
not ( w1884 , w1883 );
and ( w1885 , w15 , w1884 );
and ( w1886 , w1885 , g12 );
and ( w1887 , w1886 , w6997 );
nor ( w1888 , w1798 , w1887 );
and ( w1889 , w1888 , w1728 );
and ( w1890 , w1889 , g3 );
nor ( w1891 , w1890 , g10 );
and ( w1892 , w1891 , g12 );
and ( w1893 , w1892 , g11 );
not ( w1894 , w1795 );
and ( w1895 , w1894 , w1893 );
not ( w1896 , w1895 );
and ( w1897 , w1896 , g3 );
not ( w1898 , w663 );
and ( w1899 , w1898 , g11 );
and ( w1900 , w6161 , w1899 );
and ( w1901 , w1900 , g4 );
nor ( w1902 , w1901 , w1770 );
nor ( w1903 , w1902 , w15 );
and ( w1904 , g13 , g2 );
not ( w1905 , w1904 );
and ( w1906 , w1905 , g2 );
nor ( w1907 , w1906 , w12 );
and ( w1908 , w1907 , w1727 );
and ( w1909 , w15 , w1869 );
and ( w1910 , w1909 , w6997 );
nor ( w1911 , w1908 , w1910 );
nor ( w1912 , w1911 , g3 );
and ( w1913 , w1912 , g4 );
nor ( w1914 , w1913 , w1793 );
not ( w1915 , w1914 );
and ( w1916 , w15 , w1915 );
and ( w1917 , w1916 , w6997 );
and ( w1918 , w1917 , g12 );
and ( w1919 , w1918 , g11 );
nor ( w1920 , w1903 , w1919 );
nor ( w1921 , w1920 , g3 );
nor ( w1922 , w1921 , g3 );
nor ( w1923 , w1922 , g2 );
and ( w1924 , w1923 , w6997 );
and ( w1925 , w1924 , g12 );
and ( w1926 , w1925 , g11 );
not ( w1927 , w1897 );
and ( w1928 , w1927 , w1926 );
nor ( w1929 , w1777 , w1928 );
nor ( w1930 , w1929 , w15 );
and ( w1931 , w1930 , g12 );
and ( w1932 , w1931 , w6997 );
and ( w1933 , w1932 , g11 );
nor ( w1934 , w1773 , w1933 );
and ( w1935 , w7213 , g13 );
and ( w1936 , w1935 , w15 );
and ( w1937 , w1936 , w2606 );
nor ( w1938 , w1937 , w1733 );
and ( w1939 , w1938 , w1737 );
and ( w1940 , w1939 , g3 );
and ( w1941 , w15 , w1940 );
not ( w1942 , w1941 );
and ( w1943 , w1942 , g4 );
nor ( w1944 , w452 , w1793 );
nor ( w1945 , w1944 , g10 );
and ( w1946 , w1945 , g12 );
and ( w1947 , w1946 , g11 );
nor ( w1948 , w1943 , w1947 );
not ( w1949 , w1948 );
and ( w1950 , w1949 , g13 );
nor ( w1951 , w1950 , w1928 );
nor ( w1952 , w1951 , w12 );
and ( w1953 , w1952 , w2404 );
nor ( w1954 , w1953 , w1733 );
and ( w1955 , w1954 , w1737 );
not ( w1956 , w1955 );
and ( w1957 , w1956 , w1893 );
not ( w1958 , w1957 );
and ( w1959 , w1958 , g3 );
not ( w1960 , w1959 );
and ( w1961 , w1960 , w1926 );
not ( w1962 , w1961 );
and ( w1963 , w1934 , w1962 );
and ( w1964 , w2177 , w1963 );
not ( w1965 , w1964 );
and ( w1966 , w1965 , g4 );
nor ( w1967 , w1966 , w1772 );
not ( w1968 , w1967 );
and ( w1969 , w1968 , g2 );
and ( w1970 , w1969 , g13 );
nor ( w1971 , w1970 , w1933 );
nor ( w1972 , w1971 , w15 );
nor ( w1973 , w1935 , w1961 );
nor ( w1974 , w1973 , w12 );
and ( w1975 , w1974 , g3 );
and ( w1976 , w1975 , g4 );
not ( w1977 , w1976 );
and ( w1978 , w1977 , w15 );
nor ( w1979 , w1978 , w1728 );
nor ( w1980 , w1979 , w1887 );
not ( w1981 , w1919 );
and ( w1982 , w1980 , w1981 );
not ( w1983 , w1982 );
and ( w1984 , w1983 , w15 );
and ( w1985 , w1984 , g12 );
nor ( w1986 , w1985 , w1961 );
nor ( w1987 , w1986 , g10 );
and ( w1988 , w1987 , g11 );
nor ( w1989 , w1972 , w1988 );
not ( w1990 , w1989 );
and ( w1991 , w1990 , g12 );
and ( w1992 , w1991 , w6997 );
and ( w1993 , w1992 , g11 );
not ( w1994 , w1993 );
and ( w1995 , g13 , w1994 );
not ( w1996 , w1995 );
and ( w1997 , w1996 , g3 );
and ( w1998 , w1997 , w7213 );
and ( w1999 , w1998 , w2606 );
nor ( w2000 , w1999 , w1993 );
nor ( w2001 , w2000 , w1728 );
and ( w2002 , g2 , w7097 );
and ( w2003 , w6471 , w2002 );
and ( w2004 , w2003 , w15 );
nor ( w2005 , w2004 , w1727 );
nor ( w2006 , w2005 , w1731 );
and ( w2007 , w2006 , g10 );
and ( w2008 , w2007 , g12 );
nor ( w2009 , w2008 , w1993 );
not ( w2010 , w2009 );
and ( w2011 , w2010 , g11 );
and ( w2012 , w2011 , g4 );
and ( w2013 , w2012 , w7097 );
nor ( w2014 , w2013 , w1727 );
nor ( w2015 , w2014 , w1731 );
and ( w2016 , w2015 , g10 );
nor ( w2017 , w2016 , w1993 );
not ( w2018 , w2001 );
and ( w2019 , w2018 , w2017 );
not ( w2020 , w2019 );
and ( w2021 , w2020 , g10 );
and ( w2022 , w2021 , g12 );
nor ( w2023 , w2022 , w1993 );
not ( w2024 , w2023 );
and ( w2025 , w2024 , g11 );
and ( w2026 , w2025 , g4 );
not ( w2027 , w2026 );
and ( w2028 , w2027 , w2017 );
not ( w2029 , w2028 );
and ( w2030 , w15 , w2029 );
nor ( w2031 , w2030 , w1993 );
and ( w2032 , w452 , w7097 );
and ( w2033 , w2032 , g2 );
nor ( w2034 , w2033 , w1993 );
nor ( w2035 , w2034 , w12 );
and ( w2036 , w2035 , w3 );
and ( w2037 , w2036 , g13 );
nor ( w2038 , w2037 , w1993 );
not ( w2039 , w2038 );
and ( w2040 , w2039 , g10 );
and ( w2041 , w2040 , g12 );
nor ( w2042 , w2041 , w1993 );
not ( w2043 , w2042 );
and ( w2044 , w2043 , g11 );
not ( w2045 , w2044 );
and ( w2046 , w2031 , w2045 );
not ( w2047 , w1725 );
and ( w2048 , w2047 , w2046 );
nor ( w2049 , w2048 , w12 );
nor ( w2050 , w2049 , w1993 );
nor ( w2051 , w2050 , w1728 );
not ( w2052 , w2051 );
and ( w2053 , w2052 , w2017 );
not ( w2054 , w2053 );
and ( w2055 , w2054 , g10 );
and ( w2056 , w2055 , g12 );
nor ( w2057 , w2056 , w1993 );
not ( w2058 , w2057 );
and ( w2059 , w2058 , g11 );
nor ( w2060 , w1723 , w2059 );
nor ( w2061 , w2060 , g2 );
and ( w2062 , w2061 , w7183 );
not ( w2063 , w2062 );
and ( w2064 , w2063 , w2046 );
nor ( w2065 , w2064 , w1728 );
not ( w2066 , w2065 );
and ( w2067 , w2066 , w2017 );
not ( w2068 , w2067 );
and ( w2069 , w2068 , g10 );
and ( w2070 , w2069 , g12 );
nor ( w2071 , w2070 , w1993 );
not ( w2072 , w2071 );
and ( w2073 , w2072 , g11 );
nor ( w2074 , w1721 , w2073 );
nor ( w2075 , w2074 , g13 );
and ( w2076 , w2075 , g4 );
and ( w2077 , g10 , w2111 );
nor ( w2078 , w2077 , w1731 );
and ( w2079 , w2078 , w7102 );
and ( w2080 , w2079 , w6380 );
nor ( w2081 , w2080 , w2073 );
not ( w2082 , w2081 );
and ( w2083 , w2082 , g11 );
and ( w2084 , w2083 , w7183 );
nor ( w2085 , w2084 , w2073 );
nor ( w2086 , w2085 , g2 );
and ( w2087 , w2086 , w7097 );
and ( w2088 , w2087 , w7102 );
nor ( w2089 , w2088 , w2073 );
and ( w2090 , g8 , w5798 );
nor ( w2091 , g9 , w2090 );
nor ( w2092 , w15 , w2091 );
nor ( w2093 , w2092 , g10 );
nor ( w2094 , w2093 , w1727 );
nor ( w2095 , w2094 , w1731 );
nor ( w2096 , w2095 , w2073 );
nor ( w2097 , w2096 , g3 );
nor ( w2098 , w2097 , w370 );
nor ( w2099 , w2098 , g4 );
and ( w2100 , w2099 , w7183 );
nor ( w2101 , w2100 , w1727 );
nor ( w2102 , w2101 , w1731 );
and ( w2103 , w2102 , w6380 );
nor ( w2104 , w2103 , w2073 );
not ( w2105 , w2104 );
and ( w2106 , w2105 , g11 );
nor ( w2107 , w2106 , w1727 );
nor ( w2108 , w2107 , w1731 );
not ( w2109 , w2108 );
and ( w2110 , w2089 , w2109 );
not ( w2111 , w1727 );
and ( w2112 , w2110 , w2111 );
nor ( w2113 , w2112 , w1731 );
and ( w2114 , w2113 , w6945 );
nor ( w2115 , w2114 , w2073 );
nor ( w2116 , w2115 , g10 );
and ( w2117 , w2116 , w6471 );
nor ( w2118 , w2117 , w2073 );
and ( w2119 , w2089 , w2118 );
and ( w2120 , w6997 , w1727 );
nor ( w2121 , w2120 , w1730 );
not ( w2122 , w2121 );
and ( w2123 , w2122 , w3 );
nor ( w2124 , w2123 , w2073 );
not ( w2125 , w2124 );
and ( w2126 , w2125 , w15 );
and ( w2127 , w2126 , g4 );
and ( w2128 , w2127 , w7213 );
not ( w2129 , w2128 );
and ( w2130 , w2129 , w2089 );
nor ( w2131 , w2130 , g3 );
nor ( w2132 , w2131 , w2073 );
not ( w2133 , w2132 );
and ( w2134 , w2133 , g11 );
not ( w2135 , w2134 );
and ( w2136 , w2119 , w2135 );
nor ( w2137 , g2 , w15 );
and ( w2138 , w2091 , w7183 );
and ( w2139 , w494 , g3 );
nor ( w2140 , w2138 , w2139 );
not ( w2141 , w2137 );
and ( w2142 , w2141 , w2140 );
nor ( w2143 , w2142 , g13 );
and ( w2144 , w2143 , w7102 );
and ( w2145 , w2144 , g3 );
not ( w2146 , w2145 );
and ( w2147 , w2136 , w2146 );
not ( w2148 , w2147 );
and ( w2149 , w2148 , g10 );
not ( w2150 , w2149 );
and ( w2151 , w2150 , w2136 );
nor ( w2152 , w2151 , g4 );
and ( w2153 , w2152 , w2606 );
and ( w2154 , w2153 , w3 );
not ( w2155 , w2154 );
and ( w2156 , w2155 , w2136 );
nor ( w2157 , w2156 , g12 );
nor ( w2158 , w2157 , w2073 );
not ( w2159 , w2158 );
and ( w2160 , w2159 , g11 );
nor ( w2161 , w2076 , w2160 );
not ( w2162 , w2161 );
and ( w2163 , w2162 , w3 );
not ( w2164 , w2163 );
and ( w2165 , w2164 , w2136 );
not ( w2166 , w2165 );
and ( w2167 , w2166 , g3 );
not ( w2168 , w2167 );
and ( w2169 , w2168 , w2136 );
nor ( w2170 , w2169 , g12 );
nor ( w2171 , w2170 , w2073 );
not ( w2172 , w2171 );
and ( w2173 , w2172 , g11 );
and ( w2174 , w2173 , w15 );
and ( w2175 , w2174 , g2 );
nor ( w2176 , w2175 , w2160 );
not ( w2177 , w1729 );
and ( w2178 , w2177 , w1731 );
and ( w2179 , g10 , w3 );
and ( w2180 , w2179 , w1729 );
not ( w2181 , w2180 );
and ( w2182 , w2181 , w1731 );
nor ( w2183 , w2182 , g4 );
and ( w2184 , w2183 , w7097 );
and ( w2185 , w2184 , w7213 );
nor ( w2186 , g4 , w2185 );
nor ( w2187 , w2186 , g2 );
nor ( w2188 , w2187 , g2 );
and ( w2189 , w2188 , w7097 );
and ( w2190 , w2189 , g10 );
not ( w2191 , w2190 );
and ( w2192 , w2191 , w1729 );
not ( w2193 , w2192 );
and ( w2194 , w2193 , w1731 );
and ( w2195 , w2199 , w1729 );
not ( w2196 , w2195 );
and ( w2197 , w2196 , w1731 );
nor ( w2198 , w2178 , w2197 );
not ( w2199 , w2194 );
and ( w2200 , w2198 , w2199 );
and ( w2201 , w2200 , w1729 );
not ( w2202 , w2201 );
and ( w2203 , w2202 , w1731 );
and ( w2204 , w7183 , w1731 );
nor ( w2205 , w2204 , w150 );
nor ( w2206 , w2205 , g10 );
not ( w2207 , w2206 );
and ( w2208 , w2207 , g4 );
and ( w2209 , w2208 , w7097 );
and ( w2210 , w2209 , w7213 );
nor ( w2211 , w487 , w2210 );
and ( w2212 , w2211 , g4 );
nor ( w2213 , w2212 , g2 );
nor ( w2214 , w2213 , g2 );
and ( w2215 , w2214 , w7097 );
nor ( w2216 , w2215 , w1731 );
nor ( w2217 , w2216 , w3 );
nor ( w2218 , w2217 , w1731 );
nor ( w2219 , w2218 , w3 );
nor ( w2220 , w2219 , w2217 );
and ( w2221 , w2220 , w2357 );
nor ( w2222 , w2221 , w3 );
not ( w2223 , w2222 );
and ( w2224 , w2223 , g3 );
not ( w2225 , w2224 );
and ( w2226 , w2225 , g3 );
and ( w2227 , w2251 , g2 );
not ( w2228 , w2227 );
and ( w2229 , w2228 , g2 );
nor ( w2230 , w2229 , w2178 );
and ( w2231 , w2230 , w1729 );
not ( w2232 , w2231 );
and ( w2233 , w2232 , w1731 );
nor ( w2234 , w2233 , w2217 );
and ( w2235 , w2215 , w15 );
nor ( w2236 , w2235 , w2217 );
nor ( w2237 , w486 , g2 );
nor ( w2238 , w2237 , g2 );
and ( w2239 , w2238 , w7097 );
nor ( w2240 , w2178 , w2239 );
nor ( w2241 , w2240 , w487 );
nor ( w2242 , w2241 , g2 );
nor ( w2243 , w2242 , g2 );
and ( w2244 , w2243 , w6997 );
and ( w2245 , w2244 , w15 );
nor ( w2246 , w2229 , w2245 );
and ( w2247 , w2236 , w2246 );
and ( w2248 , w2234 , w2247 );
not ( w2249 , w2226 );
and ( w2250 , w2249 , w2248 );
not ( w2251 , w2178 );
and ( w2252 , w2251 , w2250 );
and ( w2253 , w2252 , w2248 );
and ( w2254 , w2253 , w7213 );
nor ( w2255 , w2254 , g2 );
not ( w2256 , w2255 );
and ( w2257 , w2256 , w2253 );
and ( w2258 , w1731 , w6794 );
not ( w2259 , w2258 );
and ( w2260 , w2253 , w2259 );
and ( w2261 , w2260 , w2357 );
nor ( w2262 , w2261 , w3 );
not ( w2263 , w2262 );
and ( w2264 , w2263 , w2253 );
and ( w2265 , w2257 , w2264 );
and ( w2266 , w2265 , w2357 );
nor ( w2267 , w2266 , w3 );
not ( w2268 , w2267 );
and ( w2269 , w2268 , w2253 );
and ( w2270 , w2269 , w2264 );
and ( w2271 , w2270 , w2253 );
not ( w2272 , w2203 );
and ( w2273 , w2272 , w2271 );
and ( w2274 , w2273 , w2253 );
and ( w2275 , w7094 , w2274 );
not ( w2276 , w2275 );
and ( w2277 , w2176 , w2276 );
and ( w2278 , w7183 , g3 );
not ( w2279 , w493 );
and ( w2280 , w2279 , g2 );
and ( w2281 , w2280 , w7097 );
nor ( w2282 , w2278 , w2281 );
and ( w2283 , w2282 , g4 );
and ( w2284 , w7097 , w15 );
nor ( w2285 , w2284 , w2281 );
and ( w2286 , w2285 , w7102 );
not ( w2287 , w2286 );
and ( w2288 , w2287 , g2 );
not ( w2289 , w2283 );
and ( w2290 , w2289 , w2288 );
and ( w2291 , w2290 , g13 );
nor ( w2292 , g2 , g10 );
and ( w2293 , w2292 , w7097 );
and ( w2294 , w2293 , w1727 );
nor ( w2295 , g2 , w1731 );
and ( w2296 , w2295 , w6471 );
and ( w2297 , w2296 , w15 );
nor ( w2298 , w2294 , w2297 );
not ( w2299 , w2298 );
and ( w2300 , w2299 , g4 );
and ( w2301 , w2300 , w6380 );
and ( w2302 , w2301 , w6997 );
nor ( w2303 , w2302 , w1993 );
not ( w2304 , w2303 );
and ( w2305 , w2304 , w15 );
not ( w2306 , w2305 );
and ( w2307 , w2306 , w2176 );
not ( w2308 , w2307 );
and ( w2309 , w2308 , g11 );
nor ( w2310 , w1906 , w1935 );
not ( w2311 , w2310 );
and ( w2312 , w2311 , g3 );
and ( w2313 , w1935 , w7097 );
and ( w2314 , w2313 , w2357 );
and ( w2315 , w2314 , w6997 );
nor ( w2316 , w2312 , w2315 );
not ( w2317 , w2316 );
and ( w2318 , w2317 , g4 );
and ( w2319 , w234 , w7097 );
and ( w2320 , w2319 , g2 );
and ( w2321 , w2320 , w7102 );
not ( w2322 , w2321 );
and ( w2323 , w2322 , w2176 );
and ( w2324 , w887 , w15 );
nor ( w2325 , w175 , w2324 );
not ( w2326 , w2325 );
and ( w2327 , w2326 , g2 );
and ( w2328 , w1 , w7213 );
and ( w2329 , g13 , g3 );
and ( w2330 , w2329 , w7213 );
and ( w2331 , w2330 , w7102 );
and ( w2332 , w15 , w2331 );
and ( w2333 , w2332 , w2357 );
and ( w2334 , w2333 , w6380 );
and ( w2335 , w2334 , w6997 );
and ( w2336 , w2335 , g11 );
nor ( w2337 , w2328 , w2336 );
not ( w2338 , w2337 );
and ( w2339 , w2338 , g13 );
nor ( w2340 , w2339 , w2309 );
not ( w2341 , w2340 );
and ( w2342 , w2341 , w15 );
nor ( w2343 , w2342 , w1727 );
nor ( w2344 , w2343 , w1731 );
and ( w2345 , w2344 , w6380 );
and ( w2346 , w2345 , w6997 );
nor ( w2347 , w2346 , w1993 );
and ( w2348 , w2347 , w2176 );
not ( w2349 , w2348 );
and ( w2350 , w2349 , g11 );
nor ( w2351 , w2327 , w2350 );
not ( w2352 , w2351 );
and ( w2353 , w2352 , g13 );
nor ( w2354 , w2353 , w2309 );
not ( w2355 , w2354 );
and ( w2356 , w2355 , w15 );
not ( w2357 , w1731 );
and ( w2358 , w2356 , w2357 );
and ( w2359 , w2358 , w6380 );
and ( w2360 , w2359 , w6997 );
nor ( w2361 , w2360 , w1993 );
and ( w2362 , w2361 , w2176 );
not ( w2363 , w2362 );
and ( w2364 , w2363 , g11 );
not ( w2365 , w2364 );
and ( w2366 , w2323 , w2365 );
nor ( w2367 , w2366 , w15 );
nor ( w2368 , w2367 , w2364 );
nor ( w2369 , w2368 , g10 );
not ( w2370 , w2369 );
and ( w2371 , w2370 , w2176 );
not ( w2372 , w2371 );
and ( w2373 , w2372 , g11 );
nor ( w2374 , w2318 , w2373 );
nor ( w2375 , w2374 , w15 );
nor ( w2376 , w2375 , w2364 );
nor ( w2377 , w2376 , w1731 );
and ( w2378 , w2377 , w6380 );
and ( w2379 , w2378 , w6997 );
nor ( w2380 , w2379 , w1993 );
and ( w2381 , w2380 , w2176 );
not ( w2382 , w2381 );
and ( w2383 , w2382 , g11 );
nor ( w2384 , g13 , w2383 );
not ( w2385 , w2384 );
and ( w2386 , w2385 , g3 );
and ( w2387 , w2386 , w7213 );
nor ( w2388 , w2387 , w2383 );
nor ( w2389 , w2388 , w12 );
and ( w2390 , w2389 , w2404 );
nor ( w2391 , w2390 , w2383 );
nor ( w2392 , w2391 , g12 );
and ( w2393 , w2392 , w6997 );
nor ( w2394 , w2393 , w1993 );
not ( w2395 , w2394 );
and ( w2396 , w2395 , g11 );
nor ( w2397 , w2309 , w2396 );
not ( w2398 , w2291 );
and ( w2399 , w2398 , w2397 );
not ( w2400 , w2399 );
and ( w2401 , w2400 , g2 );
nor ( w2402 , w2401 , w2396 );
nor ( w2403 , w2402 , w12 );
not ( w2404 , w1728 );
and ( w2405 , w2403 , w2404 );
nor ( w2406 , w2405 , w2383 );
nor ( w2407 , w2406 , g12 );
and ( w2408 , w2407 , w6997 );
nor ( w2409 , w2408 , w1993 );
and ( w2410 , w2409 , w2176 );
not ( w2411 , w2410 );
and ( w2412 , w2411 , g11 );
nor ( w2413 , w2412 , w2275 );
and ( w2414 , w6997 , w2413 );
and ( w2415 , w2444 , g13 );
not ( w2416 , w2415 );
and ( w2417 , w2416 , w2277 );
and ( w2418 , w2417 , w2413 );
nor ( w2419 , w2418 , w15 );
not ( w2420 , w2419 );
and ( w2421 , w2420 , w2413 );
and ( w2422 , w2421 , g3 );
nor ( w2423 , w2422 , w2414 );
and ( w2424 , w2274 , w2033 );
and ( w2425 , w2424 , w2444 );
and ( w2426 , w2425 , g13 );
not ( w2427 , w2426 );
and ( w2428 , w2427 , w2277 );
and ( w2429 , w2428 , w2413 );
nor ( w2430 , w2429 , w15 );
nor ( w2431 , w2430 , g3 );
nor ( w2432 , w2431 , w2414 );
not ( w2433 , w2432 );
and ( w2434 , w2433 , w2413 );
not ( w2435 , w2434 );
and ( w2436 , w2423 , w2435 );
and ( w2437 , w2436 , w1729 );
not ( w2438 , w2437 );
and ( w2439 , w2438 , w1731 );
not ( w2440 , w2418 );
and ( w2441 , w2440 , g3 );
not ( w2442 , w2441 );
and ( w2443 , w2442 , g3 );
not ( w2444 , w2414 );
and ( w2445 , w2444 , w2002 );
and ( w2446 , w2445 , w6471 );
not ( w2447 , w2446 );
and ( w2448 , w2447 , w2277 );
and ( w2449 , w2448 , w7097 );
nor ( w2450 , w2449 , w2414 );
and ( w2451 , w2450 , g2 );
and ( w2452 , w2413 , w7183 );
and ( w2453 , w2418 , w15 );
nor ( w2454 , w2452 , w2453 );
and ( w2455 , w2454 , w1729 );
not ( w2456 , w2455 );
and ( w2457 , w2456 , w1731 );
and ( w2458 , w2421 , w6794 );
nor ( w2459 , w2458 , w2414 );
and ( w2460 , w2468 , w2459 );
and ( w2461 , w2460 , g3 );
not ( w2462 , w2461 );
and ( w2463 , w2462 , g3 );
and ( w2464 , w2418 , w6794 );
nor ( w2465 , w2464 , w2414 );
nor ( w2466 , w2465 , g4 );
nor ( w2467 , w2466 , w2414 );
not ( w2468 , w2457 );
and ( w2469 , w2468 , w2467 );
nor ( w2470 , w2469 , g3 );
nor ( w2471 , w2470 , w2414 );
nor ( w2472 , w2471 , g4 );
nor ( w2473 , w2472 , w2414 );
not ( w2474 , w2463 );
and ( w2475 , w2474 , w2473 );
and ( w2476 , w2475 , w7213 );
not ( w2477 , w2476 );
and ( w2478 , w2477 , w2413 );
and ( w2479 , w2478 , w7102 );
nor ( w2480 , w2479 , w2414 );
nor ( w2481 , w2451 , w2480 );
nor ( w2482 , w2443 , w2481 );
nor ( w2483 , w2482 , w15 );
and ( w2484 , w2415 , g3 );
not ( w2485 , w2484 );
and ( w2486 , w2485 , w2277 );
and ( w2487 , w2486 , w2413 );
and ( w2488 , w2487 , w15 );
nor ( w2489 , w2488 , w2414 );
nor ( w2490 , w2489 , g4 );
nor ( w2491 , w2490 , w2414 );
not ( w2492 , w2483 );
and ( w2493 , w2492 , w2491 );
nor ( w2494 , w2493 , w3 );
nor ( w2495 , w2494 , w2414 );
nor ( w2496 , w2495 , g4 );
nor ( w2497 , w2496 , w2414 );
and ( w2498 , w2497 , g2 );
nor ( w2499 , w2498 , w2480 );
nor ( w2500 , w2439 , w2499 );
nor ( w2501 , w2500 , g4 );
nor ( w2502 , w2501 , w2414 );
and ( w2503 , w2502 , g2 );
nor ( w2504 , w2503 , w2480 );
nor ( w2505 , g4 , w2504 );
and ( w2506 , w2413 , w2580 );
and ( w2507 , w2588 , g13 );
not ( w2508 , w2507 );
and ( w2509 , w2508 , w2277 );
and ( w2510 , w2509 , w2413 );
and ( w2511 , w2510 , w2580 );
nor ( w2512 , w2511 , g2 );
nor ( w2513 , w2512 , g2 );
nor ( w2514 , w2513 , w2414 );
and ( w2515 , w2514 , w1729 );
not ( w2516 , w2515 );
and ( w2517 , w2516 , w1731 );
and ( w2518 , w2507 , g2 );
not ( w2519 , w2518 );
and ( w2520 , w2519 , w2277 );
and ( w2521 , w2520 , w2413 );
and ( w2522 , w2521 , w2580 );
and ( w2523 , w2522 , g2 );
nor ( w2524 , w2523 , w2504 );
nor ( w2525 , w2524 , w3 );
nor ( w2526 , w2525 , w2504 );
nor ( w2527 , w2526 , g3 );
nor ( w2528 , w2517 , w2527 );
and ( w2529 , w2528 , w2588 );
and ( w2530 , w2277 , w2580 );
and ( w2531 , w2530 , g2 );
nor ( w2532 , w2531 , w2504 );
not ( w2533 , w2532 );
and ( w2534 , w2533 , w2413 );
and ( w2535 , w2534 , w1731 );
nor ( w2536 , w2503 , w2505 );
and ( w2537 , w2536 , w6794 );
nor ( w2538 , w2535 , w2537 );
not ( w2539 , w2538 );
and ( w2540 , w2539 , w2413 );
not ( w2541 , w2540 );
and ( w2542 , w2529 , w2541 );
and ( w2543 , w2542 , w7183 );
not ( w2544 , w2522 );
and ( w2545 , w2544 , w1729 );
not ( w2546 , w2545 );
and ( w2547 , w2546 , w1731 );
and ( w2548 , w2418 , w7097 );
nor ( w2549 , w2548 , w2414 );
nor ( w2550 , w2549 , w2505 );
nor ( w2551 , w2550 , w2504 );
and ( w2552 , w2551 , w7213 );
not ( w2553 , w2552 );
and ( w2554 , w2506 , w2553 );
and ( w2555 , w2554 , w6794 );
and ( w2556 , w2555 , w7097 );
nor ( w2557 , w2556 , w2414 );
and ( w2558 , w2557 , w2588 );
not ( w2559 , w2547 );
and ( w2560 , w2559 , w2558 );
nor ( w2561 , w2560 , g3 );
nor ( w2562 , w2561 , w2504 );
and ( w2563 , w15 , w2562 );
nor ( w2564 , w2543 , w2563 );
and ( w2565 , w2564 , w7097 );
nor ( w2566 , w2565 , w2504 );
and ( w2567 , w2566 , g13 );
not ( w2568 , w2567 );
and ( w2569 , w2568 , w2277 );
and ( w2570 , w2569 , w2413 );
and ( w2571 , w2570 , w2580 );
nor ( w2572 , w2571 , g2 );
nor ( w2573 , w2572 , w2505 );
and ( w2574 , w2506 , w2573 );
nor ( w2575 , g3 , w2565 );
and ( w2576 , w2574 , w2605 );
and ( w2577 , w2576 , w6794 );
nor ( w2578 , w1731 , w2577 );
and ( w2579 , w2277 , w2602 );
not ( w2580 , w2505 );
and ( w2581 , w2579 , w2580 );
and ( w2582 , w2581 , w2413 );
and ( w2583 , w2605 , w2413 );
and ( w2584 , w2582 , w2583 );
and ( w2585 , w2584 , g2 );
and ( w2586 , w2585 , w15 );
nor ( w2587 , w2586 , w2565 );
not ( w2588 , w2504 );
and ( w2589 , w2587 , w2588 );
nor ( w2590 , w2565 , w2414 );
not ( w2591 , w2577 );
and ( w2592 , w2591 , w2590 );
and ( w2593 , w2589 , w2592 );
and ( w2594 , w2593 , g13 );
not ( w2595 , w2594 );
and ( w2596 , w2595 , w2277 );
and ( w2597 , w2596 , w2413 );
and ( w2598 , w2597 , w2506 );
nor ( w2599 , w2598 , w15 );
and ( w2600 , w2599 , w7213 );
nor ( w2601 , w2600 , w2505 );
not ( w2602 , w2578 );
and ( w2603 , w2602 , w2413 );
and ( w2604 , w2601 , w2603 );
not ( w2605 , w2575 );
and ( t_1 , w2604 , w2605 );
not ( w2606 , w12 );
and ( w2607 , w2606 , g5 );
and ( w2608 , w6997 , w2607 );
and ( w2609 , g5 , w7104 );
nor ( w2610 , g7 , w2609 );
nor ( w2611 , w2608 , w2610 );
not ( w2612 , w2611 );
and ( w2613 , g4 , w2612 );
nor ( w2614 , g10 , w2613 );
and ( w2615 , w2614 , w7183 );
and ( w2616 , g4 , w15 );
and ( w2617 , w2616 , w6997 );
and ( w2618 , w7102 , g10 );
not ( w2619 , w2610 );
and ( w2620 , w2618 , w2619 );
and ( w2621 , w2620 , w3037 );
and ( w2622 , w480 , w7213 );
nor ( w2623 , w2621 , w2622 );
nor ( w2624 , w2623 , w15 );
nor ( w2625 , w1733 , w2 );
and ( w2626 , g10 , w2625 );
nor ( w2627 , g10 , w2610 );
and ( w2628 , w2627 , w3037 );
nor ( w2629 , w2626 , w2628 );
not ( w2630 , w2629 );
and ( w2631 , w2630 , g4 );
and ( w2632 , w2629 , w7102 );
and ( w2633 , w2632 , w15 );
and ( w2634 , w2633 , w7213 );
nor ( w2635 , w2631 , w2634 );
not ( w2636 , w2635 );
and ( w2637 , w2636 , w15 );
and ( w2638 , w2637 , w7213 );
nor ( w2639 , w2624 , w2638 );
and ( w2640 , w230 , w7213 );
and ( w2641 , w2640 , w3037 );
and ( w2642 , w2641 , w15 );
and ( w2643 , w2642 , w7102 );
and ( w2644 , w2643 , g11 );
and ( w2645 , w2644 , w7097 );
not ( w2646 , w2645 );
and ( w2647 , w2646 , g10 );
not ( w2648 , w2647 );
and ( w2649 , w2648 , g10 );
and ( w2650 , w1904 , w15 );
and ( w2651 , w2650 , g11 );
and ( w2652 , w2651 , w7097 );
and ( w2653 , w2652 , w2625 );
and ( w2654 , w2653 , w6945 );
and ( w2655 , w2654 , w6997 );
and ( w2656 , w2655 , w7102 );
nor ( w2657 , w2649 , w2656 );
not ( w2658 , w2616 );
and ( w2659 , w2658 , w15 );
and ( w2660 , w2659 , g13 );
and ( w2661 , w2660 , g11 );
nor ( w2662 , w2661 , g2 );
nor ( w2663 , w2662 , g2 );
and ( w2664 , w2663 , w3037 );
not ( w2665 , w2664 );
and ( w2666 , w2665 , g10 );
not ( w2667 , w2666 );
and ( w2668 , w2667 , g10 );
nor ( w2669 , w2668 , g3 );
nor ( w2670 , w2669 , g3 );
and ( w2671 , w2657 , w2731 );
and ( w2672 , w2639 , w2671 );
nor ( w2673 , w2672 , g11 );
and ( w2674 , w2137 , g10 );
and ( w2675 , w2674 , w3037 );
and ( w2676 , w2675 , g4 );
and ( w2677 , g2 , w7183 );
and ( w2678 , w494 , w7097 );
nor ( w2679 , w2677 , w2678 );
not ( w2680 , w2679 );
and ( w2681 , w2680 , w2625 );
and ( w2682 , w2681 , g10 );
and ( w2683 , w2682 , w7102 );
and ( w2684 , w2683 , w7097 );
nor ( w2685 , w2676 , w2684 );
nor ( w2686 , w2685 , g3 );
and ( w2687 , w2686 , w7094 );
not ( w2688 , w2656 );
and ( w2689 , g11 , w2688 );
not ( w2690 , w2689 );
and ( w2691 , w2690 , w15 );
not ( w2692 , w2691 );
and ( w2693 , w2692 , w2607 );
not ( w2694 , w2693 );
and ( w2695 , w2694 , w2625 );
nor ( w2696 , w2695 , g2 );
nor ( w2697 , w2696 , g2 );
nor ( w2698 , w2697 , g10 );
nor ( w2699 , w2698 , g10 );
and ( w2700 , w2699 , g4 );
and ( w2701 , w2671 , g11 );
nor ( w2702 , w2701 , g2 );
and ( w2703 , w2702 , w6997 );
and ( w2704 , w2703 , w7097 );
nor ( w2705 , w2687 , w2704 );
nor ( w2706 , w2705 , w15 );
not ( w2707 , w2701 );
and ( w2708 , w2707 , g2 );
and ( w2709 , w2708 , w6997 );
and ( w2710 , w2709 , w15 );
and ( w2711 , w2710 , w7097 );
nor ( w2712 , w2687 , w2711 );
not ( w2713 , w2712 );
and ( w2714 , w15 , w2713 );
and ( w2715 , w2714 , w2625 );
and ( w2716 , w2708 , g10 );
and ( w2717 , w2716 , w15 );
and ( w2718 , w2717 , w3037 );
and ( w2719 , w2718 , w7097 );
nor ( w2720 , w2715 , w2719 );
nor ( w2721 , w2720 , g4 );
nor ( w2722 , w2706 , w2721 );
not ( w2723 , w2722 );
and ( w2724 , w2723 , w2625 );
nor ( w2725 , w2724 , w2719 );
nor ( w2726 , w2725 , g4 );
nor ( w2727 , w2700 , w2726 );
and ( w2728 , w2727 , w7097 );
nor ( w2729 , w2728 , g3 );
nor ( w2730 , w2687 , w2729 );
not ( w2731 , w2670 );
and ( w2732 , w2731 , w2730 );
not ( w2733 , w2673 );
and ( w2734 , w2733 , w2732 );
nor ( w2735 , w2734 , g2 );
and ( w2736 , w2735 , w7097 );
not ( w2737 , w2736 );
and ( w2738 , w2737 , w2732 );
not ( w2739 , w2613 );
and ( w2740 , w2739 , w2738 );
nor ( w2741 , w2740 , w15 );
nor ( w2742 , w2741 , w2638 );
and ( w2743 , w2742 , w2671 );
nor ( w2744 , w2743 , g11 );
not ( w2745 , w2744 );
and ( w2746 , w2745 , w2732 );
nor ( w2747 , w2746 , g2 );
and ( w2748 , w2747 , w7097 );
not ( w2749 , w2748 );
and ( w2750 , w2749 , w2732 );
not ( w2751 , w334 );
and ( w2752 , w2751 , w2750 );
not ( w2753 , w2752 );
and ( w2754 , w2753 , w2625 );
not ( w2755 , w2754 );
and ( w2756 , w2755 , w2738 );
nor ( w2757 , w2756 , w15 );
nor ( w2758 , w2757 , w2638 );
and ( w2759 , w2758 , w2671 );
nor ( w2760 , w2759 , g11 );
not ( w2761 , w2760 );
and ( w2762 , w2761 , w2732 );
nor ( w2763 , w2762 , g2 );
and ( w2764 , w2763 , w7097 );
not ( w2765 , w2764 );
and ( w2766 , w2765 , w2732 );
not ( w2767 , w2617 );
and ( w2768 , w2767 , w2766 );
not ( w2769 , w2768 );
and ( w2770 , w2769 , w2625 );
and ( w2771 , g9 , w5796 );
not ( w2772 , w2771 );
and ( w2773 , g9 , w2772 );
not ( w2774 , w2773 );
and ( w2775 , w2774 , g4 );
and ( w2776 , w2775 , w7183 );
not ( w2777 , w2776 );
and ( w2778 , w2777 , w2766 );
not ( w2779 , w2778 );
and ( w2780 , w2779 , g10 );
nor ( w2781 , w2776 , w493 );
nor ( w2782 , w2781 , g10 );
and ( w2783 , w2782 , w3037 );
nor ( w2784 , w2780 , w2783 );
nor ( w2785 , w2784 , w2607 );
not ( w2786 , w2785 );
and ( w2787 , w2786 , w2671 );
nor ( w2788 , w2787 , g11 );
not ( w2789 , w2788 );
and ( w2790 , w2789 , w2766 );
not ( w2791 , w2790 );
and ( w2792 , w2791 , g2 );
not ( w2793 , w2792 );
and ( w2794 , w2793 , w2766 );
nor ( w2795 , w2794 , g3 );
nor ( w2796 , w2770 , w2795 );
nor ( w2797 , w2796 , g11 );
not ( w2798 , w2797 );
and ( w2799 , w2798 , w2766 );
not ( w2800 , w2799 );
and ( w2801 , w2800 , g2 );
not ( w2802 , w2801 );
and ( w2803 , w2802 , w2766 );
nor ( w2804 , w2803 , g3 );
nor ( w2805 , w2615 , w2804 );
not ( w2806 , w2805 );
and ( w2807 , w2806 , w2625 );
nor ( w2808 , w2807 , w2795 );
nor ( w2809 , w2808 , g11 );
not ( w2810 , w2809 );
and ( w2811 , w2810 , w2766 );
not ( w2812 , w2811 );
and ( w2813 , w2812 , g2 );
not ( w2814 , w2813 );
and ( w2815 , w2814 , w2766 );
nor ( w2816 , w2815 , g3 );
nor ( w2817 , g3 , w2816 );
nor ( w2818 , w2817 , g11 );
nor ( w2819 , w2818 , w2816 );
not ( w2820 , w2819 );
and ( w2821 , w2820 , w2625 );
nor ( w2822 , w2821 , w2816 );
and ( w2823 , w2859 , g2 );
nor ( w2824 , w2823 , w2816 );
nor ( w2825 , w2824 , g11 );
nor ( w2826 , w2825 , w2816 );
nor ( w2827 , w2826 , w2607 );
nor ( w2828 , w2827 , w2816 );
and ( w2829 , w2828 , w6997 );
nor ( w2830 , w2829 , g10 );
nor ( w2831 , w2830 , w2816 );
and ( w2832 , w2822 , w2831 );
nor ( w2833 , w2832 , w15 );
nor ( w2834 , w2833 , w2816 );
and ( w2835 , w3031 , g2 );
not ( w2836 , w2284 );
and ( w2837 , w2836 , w15 );
and ( w2838 , w2837 , w7097 );
nor ( w2839 , w2838 , g13 );
and ( w2840 , w2839 , w3031 );
nor ( w2841 , w2840 , w2817 );
nor ( w2842 , w2841 , g2 );
nor ( w2843 , w2842 , w2817 );
and ( w2844 , w2843 , w3037 );
nor ( w2845 , w2844 , w2816 );
not ( w2846 , w2845 );
and ( w2847 , w2846 , w15 );
nor ( w2848 , w2847 , w2816 );
nor ( w2849 , w2848 , g4 );
nor ( w2850 , w2849 , w2816 );
and ( w2851 , w2850 , w6997 );
nor ( w2852 , w2851 , w2817 );
not ( w2853 , w2852 );
and ( w2854 , w2853 , g11 );
nor ( w2855 , w2835 , w2854 );
nor ( w2856 , w2855 , g10 );
and ( w2857 , w2856 , g11 );
nor ( w2858 , w2857 , g10 );
not ( w2859 , w2817 );
and ( w2860 , w2859 , w2858 );
and ( w2861 , w2860 , w15 );
and ( w2862 , w2861 , w7102 );
not ( w2863 , w2862 );
and ( w2864 , w2834 , w2863 );
and ( w2865 , w2864 , w6997 );
nor ( w2866 , w2865 , g10 );
nor ( w2867 , w2866 , w2816 );
nor ( w2868 , w2867 , g4 );
nor ( w2869 , w2868 , w2816 );
nor ( w2870 , g1 , w2817 );
and ( w2871 , w2870 , g2 );
and ( w2872 , w2871 , w7183 );
nor ( w2873 , w2872 , w2816 );
not ( w2874 , w2873 );
and ( w2875 , w2874 , w2611 );
nor ( w2876 , w2835 , w2817 );
and ( w2877 , w2876 , w7183 );
nor ( w2878 , g1 , w2816 );
nor ( w2879 , w2878 , w2817 );
and ( w2880 , w2879 , w15 );
nor ( w2881 , w2816 , w2880 );
nor ( w2882 , w2881 , g2 );
nor ( w2883 , w2882 , w2816 );
nor ( w2884 , w2883 , w2607 );
nor ( w2885 , w2884 , w2816 );
not ( w2886 , w2885 );
and ( w2887 , w2886 , g11 );
nor ( w2888 , w2887 , w2816 );
and ( w2889 , w2888 , g10 );
not ( w2890 , w2889 );
and ( w2891 , w2890 , g10 );
nor ( w2892 , w2891 , w2816 );
and ( w2893 , w2892 , w2869 );
nor ( w2894 , w2893 , g4 );
nor ( w2895 , w2894 , w2816 );
not ( w2896 , w2877 );
and ( w2897 , w2896 , w2895 );
not ( w2898 , w2897 );
and ( w2899 , w2898 , g13 );
nor ( w2900 , w2897 , g1 );
and ( w2901 , w2900 , w6471 );
nor ( w2902 , w2901 , w2816 );
not ( w2903 , w2902 );
and ( w2904 , w2903 , w2625 );
nor ( w2905 , w2904 , w2816 );
and ( w2906 , w2905 , w2895 );
not ( w2907 , w2906 );
and ( w2908 , w2907 , g11 );
nor ( w2909 , w2908 , w2816 );
not ( w2910 , w2909 );
and ( w2911 , w2910 , g10 );
nor ( w2912 , w2911 , w2816 );
and ( w2913 , w2912 , w2869 );
nor ( w2914 , w2913 , g4 );
nor ( w2915 , w2914 , w2816 );
not ( w2916 , w2899 );
and ( w2917 , w2916 , w2915 );
not ( w2918 , w2917 );
and ( w2919 , w2918 , w2625 );
nor ( w2920 , w2919 , w2816 );
and ( w2921 , w2920 , w2895 );
not ( w2922 , w2921 );
and ( w2923 , w2922 , g11 );
nor ( w2924 , w2923 , w2816 );
and ( w2925 , w2924 , g10 );
not ( w2926 , w2925 );
and ( w2927 , w2926 , g10 );
nor ( w2928 , w2927 , w2816 );
not ( w2929 , w2928 );
and ( w2930 , w2929 , w2611 );
not ( w2931 , w2930 );
and ( w2932 , w2931 , w2869 );
nor ( w2933 , w2932 , g4 );
nor ( w2934 , w2933 , w2816 );
not ( w2935 , w2875 );
and ( w2936 , w2935 , w2934 );
not ( w2937 , w2936 );
and ( w2938 , w2937 , w2625 );
nor ( w2939 , w2938 , w2816 );
and ( w2940 , w2939 , w2934 );
not ( w2941 , w2940 );
and ( w2942 , w2941 , g4 );
nor ( w2943 , w2942 , w2816 );
and ( w2944 , w2943 , w2934 );
not ( w2945 , w2944 );
and ( w2946 , w2945 , g11 );
not ( w2947 , w2946 );
and ( w2948 , w2869 , w2947 );
and ( w2949 , g11 , w2948 );
and ( w2950 , w3066 , w2625 );
and ( w2951 , w2948 , w2607 );
nor ( w2952 , w2949 , w2817 );
not ( w2953 , w2951 );
and ( w2954 , w2953 , w2952 );
and ( w2955 , w15 , w2954 );
nor ( w2956 , w2955 , w2816 );
not ( w2957 , w2956 );
and ( w2958 , w2957 , g2 );
nor ( w2959 , w2958 , w2816 );
not ( w2960 , w2959 );
and ( w2961 , w2960 , g4 );
nor ( w2962 , w2961 , g10 );
and ( w2963 , w2962 , w3031 );
nor ( w2964 , w2963 , g10 );
nor ( w2965 , w2964 , w2816 );
and ( w2966 , w2948 , w7183 );
nor ( w2967 , w2966 , w2817 );
and ( w2968 , w2967 , w3066 );
not ( w2969 , w2968 );
and ( w2970 , w2969 , w2607 );
not ( w2971 , w2970 );
and ( w2972 , w2971 , w2625 );
nor ( w2973 , w2972 , w2816 );
and ( w2974 , w2952 , w7183 );
not ( w2975 , w2948 );
and ( w2976 , w15 , w2975 );
nor ( w2977 , w2976 , w2816 );
not ( w2978 , w2974 );
and ( w2979 , w2978 , w2977 );
nor ( w2980 , w2979 , w2607 );
and ( w2981 , w2980 , g4 );
nor ( w2982 , w2981 , g10 );
nor ( w2983 , w2982 , g10 );
not ( w2984 , w2983 );
and ( w2985 , w2984 , w2869 );
and ( w2986 , w2973 , w2985 );
not ( w2987 , w2986 );
and ( w2988 , w2987 , g4 );
nor ( w2989 , w2988 , g10 );
nor ( w2990 , w2989 , g10 );
nor ( w2991 , w2990 , w2816 );
and ( w2992 , w2991 , w2869 );
and ( w2993 , w2992 , w7213 );
nor ( w2994 , w2993 , g2 );
nor ( w2995 , w2994 , w2816 );
and ( w2996 , w2965 , w2995 );
and ( w2997 , w2996 , w2869 );
not ( w2998 , w2950 );
and ( w2999 , w2998 , w2997 );
nor ( w3000 , w2999 , w2817 );
and ( w3001 , w3000 , w7183 );
not ( w3002 , w3001 );
and ( w3003 , w3002 , w2997 );
not ( w3004 , w3003 );
and ( w3005 , w3004 , g2 );
and ( w3006 , w3005 , g4 );
and ( w3007 , w3006 , w6997 );
not ( w3008 , w3007 );
and ( w3009 , w3008 , w2995 );
and ( w3010 , w3009 , w2869 );
and ( w3011 , w6997 , w3010 );
and ( w3012 , w3064 , w2952 );
and ( w3013 , w3012 , g2 );
and ( w3014 , w2948 , w3010 );
and ( w3015 , w3014 , w7213 );
nor ( w3016 , w3015 , g2 );
nor ( w3017 , w3013 , w3016 );
not ( w3018 , w3017 );
and ( w3019 , w3018 , g4 );
and ( w3020 , w3013 , w7102 );
and ( w3021 , w3014 , w7183 );
not ( w3022 , w3021 );
and ( w3023 , w3022 , w3012 );
and ( w3024 , w3023 , w3037 );
not ( w3025 , w3024 );
and ( w3026 , w3025 , w3010 );
not ( w3027 , w3020 );
and ( w3028 , w3027 , w3026 );
nor ( w3029 , w3028 , w2607 );
nor ( w3030 , w3019 , w3029 );
not ( w3031 , w2816 );
and ( w3032 , w3030 , w3031 );
and ( w3033 , w3032 , w3010 );
and ( w3034 , w3033 , w7183 );
nor ( w3035 , w3034 , w2817 );
and ( w3036 , w3035 , w3012 );
not ( w3037 , w2607 );
and ( w3038 , w3036 , w3037 );
nor ( w3039 , g10 , w3011 );
nor ( w3040 , w3038 , w3039 );
and ( w3041 , w2948 , w3040 );
and ( w3042 , w3041 , g2 );
nor ( w3043 , w3038 , w2816 );
not ( w3044 , w2625 );
and ( w3045 , w3044 , w3043 );
nor ( w3046 , w3045 , w2949 );
nor ( w3047 , w3011 , w2817 );
and ( w3048 , w3046 , w3047 );
not ( w3049 , w3042 );
and ( w3050 , w3049 , w3048 );
and ( w3051 , w3050 , w7102 );
and ( w3052 , w3043 , w3010 );
not ( w3053 , w3051 );
and ( w3054 , w3053 , w3052 );
and ( w3055 , w7102 , w3054 );
nor ( w3056 , w3055 , w3011 );
and ( w3057 , w3056 , w3046 );
and ( w3058 , w3012 , w3057 );
and ( w3059 , w3058 , g2 );
not ( w3060 , w3059 );
and ( w3061 , w3060 , w3054 );
and ( w3062 , w3061 , w15 );
nor ( w3063 , w3062 , w2817 );
not ( w3064 , w3011 );
and ( w3065 , w3063 , w3064 );
not ( w3066 , w2949 );
and ( w3067 , w3065 , w3066 );
nor ( w3068 , w3045 , w3011 );
and ( w3069 , w3067 , w3068 );
and ( t_2 , w3069 , w3056 );
nor ( w3070 , g7 , w6 );
and ( w3071 , w2609 , w6794 );
not ( w3072 , w3071 );
and ( w3073 , w3070 , w3072 );
nor ( w3074 , w3073 , w3 );
and ( w3075 , w3438 , g3 );
and ( w3076 , w6997 , w8 );
not ( w3077 , w3076 );
and ( w3078 , w3074 , w3077 );
nor ( w3079 , w3078 , g3 );
and ( w3080 , w3079 , w7213 );
nor ( w3081 , w3075 , w3080 );
and ( w3082 , w3081 , w7102 );
and ( w3083 , w3082 , w6997 );
nor ( w3084 , w3083 , g11 );
and ( w3085 , w6380 , g4 );
not ( w3086 , w3085 );
and ( w3087 , w3086 , g2 );
and ( w3088 , g12 , w7102 );
and ( w3089 , w3088 , g2 );
and ( w3090 , g12 , g4 );
and ( w3091 , w3090 , w7213 );
and ( w3092 , w3091 , g13 );
nor ( w3093 , w3089 , w3092 );
not ( w3094 , w3093 );
and ( w3095 , w3094 , g13 );
and ( w3096 , w3095 , w8 );
and ( w3097 , g12 , w6471 );
nor ( w3098 , w3097 , g4 );
not ( w3099 , w3098 );
and ( w3100 , w3099 , g3 );
nor ( w3101 , w3085 , g3 );
and ( w3102 , w3101 , g2 );
and ( w3103 , w3102 , w8 );
not ( w3104 , w3103 );
and ( w3105 , w3104 , g10 );
nor ( w3106 , g11 , g10 );
and ( w3107 , w1904 , g12 );
and ( w3108 , w3107 , g11 );
and ( w3109 , w3108 , w7102 );
and ( w3110 , w3109 , w15 );
and ( w3111 , w3107 , g1 );
and ( w3112 , w3111 , g11 );
nor ( w3113 , w3110 , w3112 );
not ( w3114 , w3113 );
and ( w3115 , w3114 , g10 );
and ( w3116 , w825 , w6997 );
and ( w3117 , w3116 , g11 );
and ( w3118 , w3117 , w7102 );
and ( w3119 , w3118 , w15 );
nor ( w3120 , w3115 , w3119 );
nor ( w3121 , w3120 , g4 );
and ( w3122 , w3121 , w15 );
and ( w3123 , w3122 , w3438 );
nor ( w3124 , w3097 , w3123 );
and ( w3125 , w3124 , g11 );
and ( w3126 , w3125 , g10 );
and ( w3127 , g13 , w6997 );
nor ( w3128 , w3127 , g10 );
and ( w3129 , w3128 , g11 );
nor ( w3130 , w3129 , w3074 );
and ( w3131 , w3130 , w15 );
not ( w3132 , w3126 );
and ( w3133 , w3132 , w3131 );
and ( w3134 , w3133 , g2 );
and ( w3135 , w3134 , w7097 );
nor ( w3136 , g13 , g2 );
and ( w3137 , w3136 , w15 );
and ( w3138 , w3137 , w7102 );
and ( w3139 , w3138 , g10 );
and ( w3140 , w3139 , w6380 );
and ( w3141 , w3140 , w7097 );
and ( w3142 , w3141 , g1 );
nor ( w3143 , w3140 , g13 );
not ( w3144 , w3143 );
and ( w3145 , w3144 , g11 );
and ( w3146 , w3145 , g10 );
and ( w3147 , w3146 , w7213 );
and ( w3148 , w3147 , w7102 );
and ( w3149 , w3148 , w15 );
and ( w3150 , w3149 , w8 );
nor ( w3151 , w3142 , w3150 );
and ( w3152 , w6471 , w3151 );
and ( w3153 , w3152 , g11 );
not ( w3154 , w3153 );
and ( w3155 , w3154 , w8 );
and ( w3156 , w3155 , w7097 );
and ( w3157 , w3156 , g10 );
and ( w3158 , w3157 , w7213 );
and ( w3159 , w3158 , w7102 );
and ( w3160 , w3159 , w15 );
nor ( w3161 , w3135 , w3160 );
nor ( w3162 , w3161 , g4 );
nor ( w3163 , g13 , w3162 );
and ( w3164 , w3163 , g11 );
and ( w3165 , w3164 , g3 );
nor ( w3166 , w824 , w3162 );
and ( w3167 , w3166 , g11 );
and ( w3168 , w3167 , w6535 );
and ( w3169 , w3168 , w3795 );
nor ( w3170 , w3169 , w3074 );
nor ( w3171 , w3170 , w3162 );
nor ( w3172 , w3090 , g2 );
nor ( w3173 , w3172 , g3 );
not ( w3174 , w3173 );
and ( w3175 , w3174 , g11 );
and ( w3176 , w3175 , w6997 );
nor ( w3177 , g13 , w3176 );
and ( w3178 , w1796 , w7213 );
and ( w3179 , w3178 , w6945 );
nor ( w3180 , w3178 , w3162 );
not ( w3181 , w3180 );
and ( w3182 , w3181 , g1 );
and ( w3183 , w3182 , w7097 );
and ( w3184 , w3183 , w3438 );
nor ( w3185 , w3184 , g10 );
and ( w3186 , w3185 , w3199 );
not ( w3187 , w3186 );
and ( w3188 , w3187 , w15 );
nor ( w3189 , w3179 , w3188 );
not ( w3190 , w3189 );
and ( w3191 , w3190 , g12 );
and ( w3192 , w3191 , w7097 );
nor ( w3193 , w3192 , g10 );
and ( w3194 , w3193 , w3199 );
not ( w3195 , w3194 );
and ( w3196 , w3195 , w15 );
and ( w3197 , w3196 , g11 );
nor ( w3198 , w3197 , g10 );
not ( w3199 , w3162 );
and ( w3200 , w3198 , w3199 );
not ( w3201 , w3177 );
and ( w3202 , w3201 , w3200 );
and ( w3203 , w3202 , g11 );
nor ( w3204 , w3203 , w3074 );
nor ( w3205 , w3204 , g10 );
not ( w3206 , w3205 );
and ( w3207 , w3206 , w15 );
nor ( w3208 , g2 , w3207 );
nor ( w3209 , w3208 , g3 );
and ( w3210 , w3209 , w3438 );
nor ( w3211 , w3210 , g10 );
not ( w3212 , w3211 );
and ( w3213 , w3212 , w15 );
not ( w3214 , w3213 );
and ( w3215 , w3171 , w3214 );
and ( w3216 , w3215 , w6997 );
nor ( w3217 , w3216 , w3074 );
and ( w3218 , w3217 , w7213 );
and ( w3219 , w3218 , g4 );
nor ( w3220 , w3219 , w3162 );
not ( w3221 , w3220 );
and ( w3222 , w3221 , w15 );
not ( w3223 , w3165 );
and ( w3224 , w3223 , w3222 );
and ( w3225 , w3224 , w6997 );
nor ( w3226 , w3225 , w3162 );
not ( w3227 , w3106 );
and ( w3228 , w3227 , w3226 );
nor ( w3229 , w3228 , g4 );
and ( w3230 , w3229 , w7213 );
and ( w3231 , w3230 , w8 );
not ( w3232 , w3231 );
and ( w3233 , w3232 , w3226 );
not ( w3234 , w3233 );
and ( w3235 , w3234 , w15 );
and ( w3236 , w3105 , w3479 );
not ( w3237 , w3236 );
and ( w3238 , w3237 , w15 );
nor ( w3239 , w3100 , w3238 );
not ( w3240 , w3239 );
and ( w3241 , w3240 , g2 );
not ( w3242 , w3097 );
and ( w3243 , w3242 , g4 );
not ( w3244 , w3243 );
and ( w3245 , w3244 , g3 );
and ( w3246 , w3097 , g4 );
and ( w3247 , w3246 , w7097 );
and ( w3248 , w3247 , w7213 );
and ( w3249 , w3248 , w8 );
not ( w3250 , w3249 );
and ( w3251 , w3250 , g10 );
and ( w3252 , w8 , g2 );
and ( w3253 , w3252 , w7102 );
nor ( w3254 , w477 , w3253 );
and ( w3255 , w555 , g12 );
and ( w3256 , w3255 , w8 );
and ( w3257 , w3256 , w6997 );
and ( w3258 , w3257 , g11 );
and ( w3259 , w3258 , w15 );
nor ( w3260 , w1796 , w3259 );
and ( w3261 , w3260 , g1 );
and ( w3262 , w3261 , g2 );
not ( w3263 , w3262 );
and ( w3264 , w3263 , w8 );
and ( w3265 , w3264 , w7097 );
and ( w3266 , w3265 , g12 );
and ( w3267 , w3266 , w6997 );
and ( w3268 , w3267 , g11 );
and ( w3269 , w3268 , w15 );
not ( w3270 , w3269 );
and ( w3271 , w3254 , w3270 );
not ( w3272 , w3271 );
and ( w3273 , w3272 , g12 );
and ( w3274 , w3273 , w6997 );
and ( w3275 , w3274 , g11 );
nor ( w3276 , w3275 , w3235 );
not ( w3277 , w3276 );
and ( w3278 , w3277 , w15 );
and ( w3279 , g12 , g2 );
nor ( w3280 , w3279 , w2 );
not ( w3281 , w3280 );
and ( w3282 , w3281 , w3 );
nor ( w3283 , w3076 , g10 );
not ( w3284 , w3282 );
and ( w3285 , w3284 , w3283 );
nor ( w3286 , w3285 , g3 );
and ( w3287 , w3286 , g13 );
nor ( w3288 , w3287 , g10 );
not ( w3289 , w3288 );
and ( w3290 , w3289 , w15 );
nor ( w3291 , w3278 , w3290 );
not ( w3292 , w3278 );
and ( w3293 , w3074 , w3292 );
not ( w3294 , w3293 );
and ( w3295 , w3294 , g3 );
and ( w3296 , w3097 , g2 );
and ( w3297 , g12 , w7213 );
and ( w3298 , w3297 , w7097 );
nor ( w3299 , w3298 , g10 );
not ( w3300 , w3299 );
and ( w3301 , w3300 , g11 );
nor ( w3302 , w3296 , w3301 );
nor ( w3303 , w3302 , g3 );
nor ( w3304 , w3303 , g10 );
not ( w3305 , w3304 );
and ( w3306 , w3305 , g11 );
nor ( w3307 , w3306 , w2 );
not ( w3308 , w3307 );
and ( w3309 , w3308 , w3 );
not ( w3310 , w3309 );
and ( w3311 , w3310 , w3283 );
nor ( w3312 , w3311 , g3 );
and ( w3313 , w3312 , g2 );
nor ( w3314 , w3301 , w2 );
not ( w3315 , w3314 );
and ( w3316 , w3315 , w3 );
not ( w3317 , w3316 );
and ( w3318 , w3317 , w3283 );
nor ( w3319 , w3318 , g3 );
and ( w3320 , w3319 , g4 );
nor ( w3321 , g2 , w3235 );
nor ( w3322 , w3321 , g12 );
nor ( w3323 , w79 , w3119 );
nor ( w3324 , w3323 , g3 );
and ( w3325 , w3324 , w3438 );
and ( w3326 , w3325 , w15 );
not ( w3327 , w3326 );
and ( w3328 , g1 , w3327 );
nor ( w3329 , w3328 , g3 );
and ( w3330 , w3329 , w3438 );
and ( w3331 , w3330 , w15 );
and ( w3332 , w3331 , g12 );
and ( w3333 , w3332 , w7213 );
nor ( w3334 , w3333 , w1904 );
and ( w3335 , w3334 , w6535 );
and ( w3336 , w3335 , w3795 );
nor ( w3337 , w3336 , w3074 );
nor ( w3338 , w3337 , w3235 );
not ( w3339 , w3338 );
and ( w3340 , w3339 , w15 );
nor ( w3341 , w3322 , w3340 );
nor ( w3342 , w3341 , w3074 );
and ( w3343 , w3342 , w6997 );
nor ( w3344 , w3343 , g10 );
not ( w3345 , w3344 );
and ( w3346 , w3345 , g11 );
and ( w3347 , w3346 , w15 );
nor ( w3348 , w3347 , w2 );
and ( w3349 , w3348 , w3795 );
nor ( w3350 , w3349 , w3074 );
nor ( w3351 , w3350 , w3278 );
nor ( w3352 , w3351 , g4 );
nor ( w3353 , w3352 , g10 );
and ( w3354 , w3353 , w3479 );
not ( w3355 , w3320 );
and ( w3356 , w3355 , w3354 );
not ( w3357 , w3356 );
and ( w3358 , w3357 , g11 );
and ( w3359 , w3358 , w15 );
nor ( w3360 , w3316 , w3278 );
not ( w3361 , w3360 );
and ( w3362 , w3361 , g4 );
not ( w3363 , w3362 );
and ( w3364 , w3363 , w3354 );
not ( w3365 , w3364 );
and ( w3366 , w3365 , w15 );
nor ( w3367 , w3359 , w3366 );
and ( w3368 , w3367 , w3354 );
not ( w3369 , w3313 );
and ( w3370 , w3369 , w3368 );
not ( w3371 , w3370 );
and ( w3372 , w3371 , g4 );
not ( w3373 , w3372 );
and ( w3374 , w3373 , w3354 );
not ( w3375 , w3374 );
and ( w3376 , w3375 , g11 );
nor ( w3377 , w3376 , w3235 );
not ( w3378 , w3377 );
and ( w3379 , w3378 , w15 );
nor ( w3380 , w3295 , w3379 );
not ( w3381 , w3380 );
and ( w3382 , w3381 , g2 );
not ( w3383 , w3382 );
and ( w3384 , w3383 , w3368 );
not ( w3385 , w3384 );
and ( w3386 , w3385 , g4 );
not ( w3387 , w3386 );
and ( w3388 , w3387 , w3354 );
not ( w3389 , w3388 );
and ( w3390 , w3389 , g11 );
and ( w3391 , w3390 , w15 );
not ( w3392 , w3391 );
and ( w3393 , w3291 , w3392 );
not ( w3394 , w3393 );
and ( w3395 , w3394 , g4 );
not ( w3396 , w3395 );
and ( w3397 , w3396 , w3354 );
not ( w3398 , w3397 );
and ( w3399 , w3398 , g11 );
nor ( w3400 , w3399 , w3235 );
nor ( w3401 , w3251 , w3400 );
and ( w3402 , w3401 , g11 );
nor ( w3403 , w3402 , w3235 );
not ( w3404 , w3403 );
and ( w3405 , w3404 , w15 );
nor ( w3406 , w3245 , w3405 );
nor ( w3407 , w3406 , g2 );
and ( w3408 , w3407 , w8 );
not ( w3409 , w3408 );
and ( w3410 , w3409 , g10 );
nor ( w3411 , w3410 , w3400 );
and ( w3412 , w3411 , g11 );
nor ( w3413 , w3412 , w3235 );
not ( w3414 , w3413 );
and ( w3415 , w3414 , w15 );
nor ( w3416 , w3241 , w3415 );
not ( w3417 , w3416 );
and ( w3418 , w3417 , w8 );
not ( w3419 , w3418 );
and ( w3420 , w3419 , g10 );
nor ( w3421 , w3420 , w3400 );
and ( w3422 , w3421 , g11 );
and ( w3423 , w3422 , w15 );
nor ( w3424 , w3096 , w3423 );
not ( w3425 , w3424 );
and ( w3426 , w3425 , g3 );
and ( w3427 , g12 , w6535 );
and ( w3428 , w3427 , w3795 );
nor ( w3429 , w3428 , w3074 );
not ( w3430 , w3423 );
and ( w3431 , w3430 , g10 );
nor ( w3432 , w3431 , w3400 );
nor ( w3433 , w3429 , w3432 );
not ( w3434 , w3433 );
and ( w3435 , w3434 , g13 );
nor ( w3436 , w578 , w78 );
nor ( w3437 , w3436 , g13 );
not ( w3438 , w3074 );
and ( w3439 , w3437 , w3438 );
nor ( w3440 , w3439 , w3238 );
not ( w3441 , w3440 );
and ( w3442 , w3441 , g2 );
and ( w3443 , w3442 , g4 );
and ( w3444 , w3443 , w7097 );
not ( w3445 , w3444 );
and ( w3446 , w3445 , g10 );
and ( w3447 , w3446 , w3479 );
not ( w3448 , w3447 );
and ( w3449 , w3448 , w15 );
nor ( w3450 , w3435 , w3449 );
not ( w3451 , w3450 );
and ( w3452 , w3451 , g2 );
and ( w3453 , g12 , w7097 );
and ( w3454 , w887 , w7213 );
and ( w3455 , w3453 , w3454 );
and ( w3456 , w3455 , g13 );
and ( w3457 , w3456 , w8 );
nor ( w3458 , w3457 , w3423 );
and ( w3459 , w3458 , w6794 );
nor ( w3460 , w3459 , g2 );
and ( w3461 , w3460 , g4 );
and ( w3462 , w79 , w7213 );
and ( w3463 , w3462 , w7097 );
not ( w3464 , w3463 );
and ( w3465 , w3464 , g10 );
not ( w3466 , w3465 );
and ( w3467 , w3466 , w15 );
nor ( w3468 , w3279 , w3467 );
and ( w3469 , w3468 , w6535 );
and ( w3470 , w3469 , w3795 );
nor ( w3471 , w3470 , w3074 );
and ( w3472 , w4133 , g10 );
not ( w3473 , w3471 );
and ( w3474 , w3473 , w3472 );
nor ( w3475 , w3474 , g4 );
and ( w3476 , w3475 , w7097 );
not ( w3477 , w3476 );
and ( w3478 , w3477 , g10 );
not ( w3479 , w3235 );
and ( w3480 , w3478 , w3479 );
not ( w3481 , w3480 );
and ( w3482 , w3481 , w15 );
nor ( w3483 , w3461 , w3482 );
nor ( w3484 , w3483 , g3 );
not ( w3485 , w3484 );
and ( w3486 , w3485 , g10 );
nor ( w3487 , w3486 , w3400 );
and ( w3488 , w3487 , w15 );
nor ( w3489 , w3452 , w3488 );
not ( w3490 , w3489 );
and ( w3491 , w3490 , g4 );
nor ( w3492 , w3491 , w3482 );
nor ( w3493 , w3492 , g3 );
not ( w3494 , w3493 );
and ( w3495 , w3494 , g10 );
nor ( w3496 , w3495 , w3400 );
and ( w3497 , w3496 , g11 );
and ( w3498 , w3497 , w15 );
nor ( w3499 , w3426 , w3498 );
and ( w3500 , w3499 , g10 );
nor ( w3501 , w3500 , w3400 );
and ( w3502 , w3501 , g11 );
and ( w3503 , w3502 , w15 );
not ( w3504 , w3503 );
and ( w3505 , w3504 , g10 );
nor ( w3506 , w3505 , w3400 );
nor ( w3507 , w3506 , g12 );
nor ( w3508 , w3507 , g13 );
and ( w3509 , w3508 , w7213 );
nor ( w3510 , w3509 , w2 );
and ( w3511 , w3510 , w3795 );
nor ( w3512 , w3511 , w3074 );
nor ( w3513 , w3512 , w3503 );
not ( w3514 , w3513 );
and ( w3515 , w3514 , g3 );
nor ( w3516 , w3515 , w3498 );
and ( w3517 , w3516 , g10 );
nor ( w3518 , w3517 , w3400 );
and ( w3519 , w3518 , g11 );
nor ( w3520 , w3519 , w3235 );
not ( w3521 , w3520 );
and ( w3522 , w3521 , w15 );
nor ( w3523 , w824 , w3522 );
nor ( w3524 , w3523 , g2 );
nor ( w3525 , w3524 , w2 );
and ( w3526 , w3525 , w3795 );
nor ( w3527 , w3526 , w3074 );
nor ( w3528 , w3527 , w3503 );
not ( w3529 , w3528 );
and ( w3530 , w3529 , g3 );
nor ( w3531 , w3530 , w3498 );
and ( w3532 , w3531 , g10 );
nor ( w3533 , w3532 , w3400 );
and ( w3534 , w3533 , g11 );
nor ( w3535 , w3534 , w3235 );
not ( w3536 , w3535 );
and ( w3537 , w3536 , w15 );
nor ( w3538 , w3087 , w3537 );
and ( w3539 , w3538 , w6535 );
and ( w3540 , w3539 , w3795 );
nor ( w3541 , w3540 , w3074 );
nor ( w3542 , w3541 , w3503 );
not ( w3543 , w3542 );
and ( w3544 , w3543 , g3 );
nor ( w3545 , w3544 , w3498 );
and ( w3546 , w3545 , g10 );
nor ( w3547 , w3546 , w3400 );
and ( w3548 , w3547 , g11 );
nor ( w3549 , w3548 , w3235 );
not ( w3550 , w3549 );
and ( w3551 , w3550 , w15 );
nor ( w3552 , w3084 , w3551 );
not ( w3553 , w3552 );
and ( w3554 , w3553 , w15 );
not ( w3555 , w201 );
and ( w3556 , w3555 , w3554 );
nor ( w3557 , w3556 , g2 );
and ( w3558 , w3557 , w6997 );
nor ( w3559 , w3558 , g11 );
nor ( w3560 , w3559 , w3551 );
not ( w3561 , w3560 );
and ( w3562 , w3561 , w15 );
nor ( w3563 , w3562 , g12 );
nor ( w3564 , w3562 , g8 );
and ( w3565 , w3564 , w5798 );
nor ( w3566 , w3563 , w3565 );
nor ( w3567 , w3566 , g2 );
nor ( w3568 , w3567 , w3565 );
not ( w3569 , w3568 );
and ( w3570 , w3569 , g10 );
and ( w3571 , w3567 , w6997 );
and ( w3572 , w3571 , w6535 );
nor ( w3573 , w3572 , w3565 );
nor ( w3574 , w3573 , w8 );
nor ( w3575 , w3574 , w3565 );
not ( w3576 , w3575 );
and ( w3577 , w3576 , g4 );
nor ( w3578 , w3570 , w3577 );
not ( w3579 , w3578 );
and ( w3580 , w3579 , g3 );
nor ( w3581 , w3580 , w3565 );
nor ( w3582 , w3566 , g3 );
and ( w3583 , w3582 , w6997 );
and ( w3584 , w3603 , g2 );
nor ( w3585 , w3584 , w3565 );
not ( w3586 , w3585 );
and ( w3587 , w3586 , w3074 );
and ( w3588 , w3587 , g10 );
nor ( w3589 , w3588 , w3565 );
not ( w3590 , w3589 );
and ( w3591 , w3590 , g3 );
nor ( w3592 , w3591 , w3565 );
nor ( w3593 , w3566 , g10 );
nor ( w3594 , w3565 , w3593 );
nor ( w3595 , w3594 , g3 );
nor ( w3596 , w3595 , w3565 );
not ( w3597 , w3596 );
and ( w3598 , w3597 , w3074 );
nor ( w3599 , w3598 , w3565 );
not ( w3600 , w3599 );
and ( w3601 , w3600 , g4 );
nor ( w3602 , w3601 , w3565 );
not ( w3603 , w3566 );
and ( w3604 , w3603 , g3 );
nor ( w3605 , w3604 , w3565 );
not ( w3606 , w3605 );
and ( w3607 , w3606 , g2 );
nor ( w3608 , w3582 , w3565 );
nor ( w3609 , w3608 , g4 );
nor ( w3610 , w3609 , w3565 );
nor ( w3611 , w3565 , w78 );
nor ( w3612 , w3611 , w3562 );
and ( w3613 , w3612 , w7213 );
nor ( w3614 , w3613 , w3565 );
not ( w3615 , w3614 );
and ( w3616 , w3615 , g10 );
nor ( w3617 , w3616 , w3565 );
nor ( w3618 , w3614 , g10 );
nor ( w3619 , w3618 , w3565 );
nor ( w3620 , w3619 , g4 );
nor ( w3621 , w3620 , w3565 );
not ( w3622 , w3621 );
and ( w3623 , w3622 , g3 );
nor ( w3624 , w3623 , w3565 );
and ( w3625 , w4777 , g12 );
not ( w3626 , w3625 );
and ( w3627 , g12 , w3626 );
and ( w3628 , w3627 , w3659 );
nor ( w3629 , w3628 , w3565 );
nor ( w3630 , w3629 , g2 );
nor ( w3631 , w3630 , w3565 );
and ( w3632 , w3641 , g10 );
nor ( w3633 , w3632 , w3565 );
and ( w3634 , w3612 , g2 );
nor ( w3635 , w3634 , w3565 );
nor ( w3636 , w3635 , g10 );
nor ( w3637 , w3636 , w3565 );
not ( w3638 , w3637 );
and ( w3639 , w3638 , g4 );
nor ( w3640 , w3639 , w3565 );
not ( w3641 , w3631 );
and ( w3642 , w3641 , g3 );
nor ( w3643 , w3642 , w3565 );
not ( w3644 , w3629 );
and ( w3645 , w3644 , g2 );
and ( w3646 , w3645 , w7097 );
nor ( w3647 , w3646 , w3565 );
not ( w3648 , w3647 );
and ( w3649 , w3648 , g4 );
nor ( w3650 , w3649 , w3565 );
and ( w3651 , w3643 , w3650 );
not ( w3652 , w3651 );
and ( w3653 , w3652 , g4 );
nor ( w3654 , w3653 , w3565 );
nor ( w3655 , g1 , w3625 );
nor ( w3656 , w3655 , w3565 );
nor ( w3657 , w3656 , w3562 );
and ( w3658 , w3657 , g3 );
not ( w3659 , w3562 );
and ( w3660 , w78 , w3659 );
nor ( w3661 , w3660 , g10 );
nor ( w3662 , w3661 , g10 );
and ( w3663 , w3563 , w7183 );
and ( w3664 , w3663 , g10 );
nor ( w3665 , w3662 , w3664 );
not ( w3666 , w3665 );
and ( w3667 , w3666 , g3 );
nor ( w3668 , w3436 , g10 );
not ( w3669 , w3668 );
and ( w3670 , w3669 , w8 );
not ( w3671 , w3670 );
and ( w3672 , w3671 , w3074 );
nor ( w3673 , w3664 , w3672 );
and ( w3674 , g12 , w8 );
nor ( w3675 , w3674 , g10 );
not ( w3676 , w3675 );
and ( w3677 , w3673 , w3676 );
nor ( w3678 , w3677 , w3562 );
and ( w3679 , w3678 , w7097 );
and ( w3680 , w3679 , w7102 );
not ( w3681 , w3680 );
and ( w3682 , w3681 , w8 );
not ( w3683 , w3682 );
and ( w3684 , w3683 , w3074 );
and ( w3685 , w3684 , w7213 );
nor ( w3686 , w3667 , w3685 );
nor ( w3687 , w3686 , g4 );
not ( w3688 , w3687 );
and ( w3689 , w3688 , w8 );
not ( w3690 , w3689 );
and ( w3691 , w3690 , w3074 );
and ( w3692 , w3691 , g11 );
and ( w3693 , w3692 , w7213 );
nor ( w3694 , w3693 , w3565 );
not ( w3695 , w3658 );
and ( w3696 , w3695 , w3694 );
not ( w3697 , w3696 );
and ( w3698 , w3697 , g2 );
and ( w3699 , w3698 , w7102 );
nor ( w3700 , w3699 , w3565 );
and ( w3701 , w3700 , w3694 );
not ( w3702 , w3701 );
and ( w3703 , w3702 , g11 );
not ( w3704 , w3703 );
and ( w3705 , w3654 , w3704 );
not ( w3706 , w3705 );
and ( w3707 , w3706 , g10 );
nor ( w3708 , w3707 , w3565 );
and ( w3709 , w3657 , w7097 );
nor ( w3710 , w3709 , w3565 );
nor ( w3711 , w3710 , g10 );
nor ( w3712 , w3711 , w3565 );
not ( w3713 , w3712 );
and ( w3714 , w3713 , g2 );
and ( w3715 , w3714 , w7102 );
nor ( w3716 , w3715 , w3565 );
and ( w3717 , w3716 , w8 );
not ( w3718 , w3717 );
and ( w3719 , w3718 , w3074 );
nor ( w3720 , w3719 , w3565 );
and ( w3721 , w3720 , w3831 );
not ( w3722 , w3721 );
and ( w3723 , w3722 , g11 );
nor ( w3724 , w3723 , g10 );
nor ( w3725 , w3724 , g10 );
nor ( w3726 , w3725 , w3565 );
and ( w3727 , w3708 , w3726 );
and ( w3728 , w3727 , w8 );
not ( w3729 , w3728 );
and ( w3730 , w3729 , w3074 );
nor ( w3731 , w3730 , w3565 );
not ( w3732 , w3731 );
and ( w3733 , w3732 , g11 );
and ( w3734 , w3640 , w3739 );
nor ( w3735 , w3734 , g3 );
nor ( w3736 , w3735 , w3565 );
nor ( w3737 , w3736 , w8 );
nor ( w3738 , w3737 , w3565 );
not ( w3739 , w3733 );
and ( w3740 , w3738 , w3739 );
not ( w3741 , w3740 );
and ( w3742 , w3741 , g11 );
not ( w3743 , w3742 );
and ( w3744 , w3633 , w3743 );
not ( w3745 , w3744 );
and ( w3746 , w3745 , g4 );
nor ( w3747 , w3746 , w3733 );
nor ( w3748 , w3747 , g3 );
nor ( w3749 , w3748 , w3565 );
nor ( w3750 , w3749 , w8 );
nor ( w3751 , w3750 , w3733 );
not ( w3752 , w3751 );
and ( w3753 , w3752 , g11 );
and ( w3754 , w3624 , w3767 );
nor ( w3755 , w3754 , w8 );
nor ( w3756 , w3755 , w3733 );
not ( w3757 , w3756 );
and ( w3758 , w3757 , g11 );
not ( w3759 , w3758 );
and ( w3760 , w3617 , w3759 );
not ( w3761 , w3760 );
and ( w3762 , w3761 , g4 );
nor ( w3763 , w3762 , w3758 );
not ( w3764 , w3763 );
and ( w3765 , w3764 , g3 );
nor ( w3766 , w3765 , w3565 );
not ( w3767 , w3753 );
and ( w3768 , w3766 , w3767 );
nor ( w3769 , w3768 , w8 );
nor ( w3770 , w3769 , w3733 );
not ( w3771 , w3770 );
and ( w3772 , w3771 , g11 );
and ( w3773 , w3610 , w3814 );
not ( w3774 , w3773 );
and ( w3775 , w3774 , g11 );
and ( w3776 , w3775 , g10 );
nor ( w3777 , w3776 , w3565 );
nor ( w3778 , w3777 , w8 );
nor ( w3779 , w3778 , w3693 );
nor ( w3780 , w3779 , g4 );
nor ( w3781 , w3780 , w3772 );
nor ( w3782 , w3781 , g2 );
and ( w3783 , w3782 , g10 );
nor ( w3784 , w3783 , w3565 );
and ( w3785 , w3563 , w6535 );
nor ( w3786 , w3785 , w3565 );
nor ( w3787 , w3786 , w8 );
nor ( w3788 , w3787 , w3565 );
not ( w3789 , w3788 );
and ( w3790 , w3789 , g3 );
nor ( w3791 , w3790 , w3565 );
and ( w3792 , w3584 , w886 );
nor ( w3793 , w3792 , w3772 );
nor ( w3794 , w3793 , w2 );
not ( w3795 , w8 );
and ( w3796 , w3794 , w3795 );
not ( w3797 , w3796 );
and ( w3798 , w3797 , w3694 );
nor ( w3799 , w3798 , g3 );
nor ( w3800 , w3799 , w3565 );
nor ( w3801 , w3800 , g10 );
nor ( w3802 , w3801 , w3565 );
nor ( w3803 , w3802 , g4 );
nor ( w3804 , w3803 , w3565 );
and ( w3805 , w3804 , w3814 );
not ( w3806 , w3805 );
and ( w3807 , w3806 , g11 );
not ( w3808 , w3807 );
and ( w3809 , w3791 , w3808 );
nor ( w3810 , w3809 , g10 );
nor ( w3811 , w3810 , w3565 );
nor ( w3812 , w3811 , g4 );
nor ( w3813 , w3812 , w3565 );
not ( w3814 , w3772 );
and ( w3815 , w3813 , w3814 );
not ( w3816 , w3815 );
and ( w3817 , w3816 , g11 );
and ( w3818 , w3784 , w3844 );
not ( w3819 , w3607 );
and ( w3820 , w3819 , w3818 );
nor ( w3821 , w3820 , w8 );
nor ( w3822 , w3587 , w3693 );
not ( w3823 , w3565 );
and ( w3824 , w3822 , w3823 );
nor ( w3825 , w3824 , g4 );
nor ( w3826 , w3825 , w3565 );
not ( w3827 , w3826 );
and ( w3828 , w3827 , g11 );
and ( w3829 , w3828 , w7097 );
nor ( w3830 , w3829 , w3565 );
not ( w3831 , w3693 );
and ( w3832 , w3830 , w3831 );
not ( w3833 , w3832 );
and ( w3834 , w3833 , g10 );
nor ( w3835 , w3834 , w3565 );
and ( w3836 , w3835 , w3844 );
not ( w3837 , w3821 );
and ( w3838 , w3837 , w3836 );
not ( w3839 , w3838 );
and ( w3840 , w3839 , g10 );
nor ( w3841 , w3840 , w3565 );
nor ( w3842 , w3841 , g4 );
nor ( w3843 , w3842 , w3565 );
not ( w3844 , w3817 );
and ( w3845 , w3843 , w3844 );
not ( w3846 , w3845 );
and ( w3847 , w3846 , g11 );
and ( w3848 , w3602 , w3866 );
not ( w3849 , w3848 );
and ( w3850 , w3849 , g11 );
not ( w3851 , w3850 );
and ( w3852 , w3592 , w3851 );
not ( w3853 , w3852 );
and ( w3854 , w3853 , g4 );
nor ( w3855 , w3854 , w3847 );
not ( w3856 , w3855 );
and ( w3857 , w3856 , g11 );
nor ( w3858 , w3583 , w3857 );
nor ( w3859 , w3858 , w2 );
nor ( w3860 , w3859 , w3565 );
nor ( w3861 , w3860 , w8 );
nor ( w3862 , w3861 , w3857 );
not ( w3863 , w3862 );
and ( w3864 , w3863 , g4 );
nor ( w3865 , w3864 , w3565 );
not ( w3866 , w3847 );
and ( w3867 , w3865 , w3866 );
not ( w3868 , w3867 );
and ( w3869 , w3868 , g11 );
not ( w3870 , w3869 );
and ( w3871 , w3581 , w3870 );
nor ( w3872 , w3871 , w2 );
nor ( w3873 , w3872 , w3565 );
nor ( w3874 , w3873 , w8 );
nor ( w3875 , w3874 , w3857 );
not ( w3876 , w3875 );
and ( w3877 , w3876 , g4 );
nor ( w3878 , w3877 , w3847 );
not ( w3879 , w3878 );
and ( t_3 , w3879 , g11 );
and ( w3880 , g12 , w15 );
not ( w3881 , w3880 );
and ( w3882 , w15 , w3881 );
and ( w3883 , w3882 , g2 );
nor ( w3884 , g12 , g2 );
and ( w3885 , g4 , w7213 );
and ( w3886 , w3884 , w3885 );
nor ( w3887 , w3883 , w3886 );
not ( w3888 , w3887 );
and ( w3889 , w3888 , g10 );
and ( w3890 , w3886 , w6997 );
and ( w3891 , w1904 , w7183 );
and ( w3892 , w3891 , g4 );
and ( w3893 , w3892 , w6945 );
and ( w3894 , w3893 , w7097 );
and ( w3895 , w650 , g2 );
and ( w3896 , w3895 , w7097 );
and ( w3897 , w3896 , w7102 );
and ( w3898 , w3897 , w7183 );
and ( w3899 , w160 , g4 );
and ( w3900 , w3899 , w7097 );
and ( w3901 , w3900 , w6997 );
and ( w3902 , w3901 , g11 );
and ( w3903 , w3902 , w8 );
and ( w3904 , w3903 , g13 );
and ( w3905 , w3453 , w6945 );
and ( w3906 , w3905 , w6471 );
and ( w3907 , w3906 , w15 );
and ( w3908 , w3907 , w8 );
nor ( w3909 , w3908 , w2324 );
nor ( w3910 , w3909 , g1 );
and ( w3911 , w3910 , w6471 );
and ( w3912 , w3911 , g4 );
and ( w3913 , w3912 , w6997 );
and ( w3914 , w3913 , g11 );
and ( w3915 , w3914 , w8 );
nor ( w3916 , w3904 , w3915 );
not ( w3917 , w3916 );
and ( w3918 , w3917 , w15 );
nor ( w3919 , w3898 , w3918 );
nor ( w3920 , w3919 , g10 );
and ( w3921 , w3920 , g11 );
and ( w3922 , w3921 , w8 );
nor ( w3923 , w3894 , w3922 );
not ( w3924 , w3923 );
and ( w3925 , w3924 , g10 );
nor ( w3926 , w3925 , w3922 );
not ( w3927 , w3926 );
and ( w3928 , w3927 , g11 );
and ( w3929 , w3928 , w8 );
nor ( w3930 , w3890 , w3929 );
nor ( w3931 , w3930 , w15 );
and ( w3932 , w3931 , w6997 );
nor ( w3933 , w3932 , w3929 );
and ( w3934 , w4553 , g4 );
nor ( w3935 , w3934 , g10 );
nor ( w3936 , w3935 , w3929 );
nor ( w3937 , w3929 , g4 );
nor ( w3938 , w3936 , w3937 );
and ( w3939 , w3938 , g3 );
not ( w3940 , w3939 );
and ( w3941 , w3940 , g3 );
and ( w3942 , w3941 , g12 );
and ( w3943 , w3942 , w15 );
not ( w3944 , w3943 );
and ( w3945 , g12 , w3944 );
and ( w3946 , w3945 , g3 );
nor ( w3947 , g4 , w493 );
nor ( w3948 , w3947 , w3929 );
and ( w3949 , w3948 , w7213 );
not ( w3950 , w228 );
and ( w3951 , w3949 , w3950 );
not ( w3952 , w3951 );
and ( w3953 , w3952 , w2625 );
nor ( w3954 , w3953 , w3929 );
and ( w3955 , w3954 , w6997 );
and ( w3956 , w3955 , w7213 );
nor ( w3957 , w452 , w3956 );
and ( w3958 , w3957 , w7097 );
and ( w3959 , w3958 , w6997 );
and ( w3960 , w3959 , w2625 );
nor ( w3961 , w3960 , w3929 );
and ( w3962 , w3961 , w7213 );
not ( w3963 , w3962 );
and ( w3964 , w3963 , g4 );
and ( w3965 , w829 , w2625 );
and ( w3966 , w3965 , w15 );
and ( w3967 , w3966 , w7097 );
and ( w3968 , w3967 , g10 );
and ( w3969 , w829 , g3 );
and ( w3970 , w3969 , w7183 );
and ( w3971 , w3970 , w2625 );
and ( w3972 , w3971 , w6997 );
nor ( w3973 , w3972 , w3929 );
not ( w3974 , w3968 );
and ( w3975 , w3974 , w3973 );
nor ( w3976 , w3975 , g4 );
nor ( w3977 , w3976 , w3929 );
not ( w3978 , w3964 );
and ( w3979 , w3978 , w3977 );
not ( w3980 , w3979 );
and ( w3981 , w3980 , w2625 );
and ( w3982 , w1747 , g10 );
nor ( w3983 , w3982 , w3929 );
nor ( w3984 , w3983 , g3 );
nor ( w3985 , w3984 , g3 );
and ( w3986 , w3985 , g12 );
and ( w3987 , w3986 , w15 );
not ( w3988 , w3981 );
and ( w3989 , w3988 , w3987 );
not ( w3990 , w3989 );
and ( w3991 , w3990 , g10 );
nor ( w3992 , w3991 , w3929 );
nor ( w3993 , w3992 , g3 );
nor ( w3994 , w3993 , g3 );
and ( w3995 , w3994 , g12 );
and ( w3996 , w3995 , w15 );
not ( w3997 , w3996 );
and ( w3998 , g2 , w3997 );
and ( w3999 , w3998 , w7097 );
nor ( w4000 , w3886 , w3929 );
not ( w4001 , w4000 );
and ( w4002 , w4001 , w2625 );
nor ( w4003 , w4002 , w3929 );
not ( w4004 , w4003 );
and ( w4005 , w4004 , w15 );
and ( w4006 , w4005 , w7097 );
and ( w4007 , w4006 , w6997 );
nor ( w4008 , w4007 , w3929 );
not ( w4009 , w93 );
and ( w4010 , w4009 , w4008 );
nor ( w4011 , w4010 , g12 );
nor ( w4012 , w4011 , w3929 );
not ( w4013 , w4012 );
and ( w4014 , w4013 , w2625 );
nor ( w4015 , w4014 , w3929 );
nor ( w4016 , w4015 , g3 );
and ( w4017 , w4016 , w6997 );
nor ( w4018 , w4017 , w3929 );
not ( w4019 , w3999 );
and ( w4020 , w4019 , w4018 );
not ( w4021 , w4020 );
and ( w4022 , w4021 , g4 );
and ( w4023 , w4022 , w6997 );
nor ( w4024 , w3946 , w4023 );
not ( w4025 , w4024 );
and ( w4026 , w4025 , w2625 );
and ( w4027 , g3 , w6380 );
and ( w4028 , w4027 , w8 );
nor ( w4029 , w4028 , w3929 );
not ( w4030 , w4029 );
and ( w4031 , w4030 , g4 );
nor ( w4032 , w367 , w3929 );
not ( w4033 , w4032 );
and ( w4034 , w4033 , w2625 );
not ( w4035 , w370 );
and ( w4036 , w4035 , w8 );
and ( w4037 , w4036 , w7102 );
and ( w4038 , w4037 , w5796 );
and ( w4039 , w4038 , w15 );
nor ( w4040 , w4034 , w4039 );
nor ( w4041 , w4040 , g12 );
not ( w4042 , w4041 );
and ( w4043 , w4042 , w3937 );
nor ( w4044 , w4043 , g4 );
and ( w4045 , w4044 , w6997 );
and ( w4046 , w4045 , w5796 );
and ( w4047 , w4046 , w15 );
nor ( w4048 , w4047 , w3929 );
not ( w4049 , w4031 );
and ( w4050 , w4049 , w4048 );
nor ( w4051 , w4050 , g10 );
and ( w4052 , w4051 , w5796 );
and ( w4053 , w4052 , w15 );
nor ( w4054 , w4053 , w3929 );
not ( w4055 , w4026 );
and ( w4056 , w4055 , w4054 );
not ( w4057 , w4056 );
and ( w4058 , w4057 , g4 );
not ( w4059 , w4058 );
and ( w4060 , w4059 , w4048 );
nor ( w4061 , w4060 , g10 );
and ( w4062 , w4061 , w5796 );
and ( w4063 , w4062 , w15 );
nor ( w4064 , w4063 , w3929 );
and ( w4065 , w3933 , w4064 );
not ( w4066 , w4065 );
and ( w4067 , w4066 , g4 );
nor ( w4068 , w829 , w3929 );
not ( w4069 , w4068 );
and ( w4070 , w4069 , g10 );
and ( w4071 , w3884 , w6997 );
and ( w4072 , w4071 , w7102 );
and ( w4073 , w4072 , g3 );
and ( w4074 , w4073 , w2625 );
nor ( w4075 , w4070 , w4074 );
nor ( w4076 , w4075 , w15 );
and ( w4077 , w4076 , w7102 );
and ( w4078 , w2625 , w7213 );
and ( w4079 , w4078 , g3 );
and ( w4080 , w4079 , w7102 );
and ( w4081 , w4080 , w5796 );
and ( w4082 , w4081 , w15 );
nor ( w4083 , w3252 , w4082 );
and ( w4084 , w4083 , w6380 );
and ( w4085 , w4553 , g12 );
not ( w4086 , w4085 );
and ( w4087 , w4086 , g3 );
and ( w4088 , w4087 , g10 );
not ( w4089 , w4084 );
and ( w4090 , w4089 , w4088 );
and ( w4091 , w3977 , w6380 );
nor ( w4092 , w4091 , w3996 );
and ( w4093 , w4092 , w7097 );
not ( w4094 , w4093 );
and ( w4095 , w4094 , w4064 );
not ( w4096 , w4095 );
and ( w4097 , w4096 , w15 );
nor ( w4098 , w4097 , w3929 );
not ( w4099 , w4090 );
and ( w4100 , w4099 , w4098 );
nor ( w4101 , w4100 , g4 );
not ( w4102 , w4101 );
and ( w4103 , w4102 , w3977 );
not ( w4104 , w4103 );
and ( w4105 , w4104 , g10 );
not ( w4106 , w4105 );
and ( w4107 , w4106 , w4064 );
nor ( w4108 , w4107 , g8 );
and ( w4109 , w4108 , w15 );
nor ( w4110 , w4109 , w3929 );
not ( w4111 , w4077 );
and ( w4112 , w4111 , w4110 );
and ( w4113 , w4112 , w3977 );
not ( w4114 , w4113 );
and ( w4115 , w4114 , g3 );
and ( w4116 , w8 , w3885 );
and ( w4117 , w4116 , g10 );
nor ( w4118 , w3252 , w4117 );
not ( w4119 , w150 );
and ( w4120 , w4119 , g10 );
not ( w4121 , w4120 );
and ( w4122 , w2295 , w4121 );
and ( w4123 , w4122 , w3885 );
nor ( w4124 , w4120 , g3 );
and ( w4125 , w4123 , w4124 );
nor ( w4126 , w4125 , g12 );
nor ( w4127 , w4126 , g3 );
and ( w4128 , w4127 , g4 );
and ( w4129 , w4128 , g10 );
and ( w4130 , w4129 , w5796 );
and ( w4131 , w4130 , w15 );
nor ( w4132 , w4131 , w3929 );
not ( w4133 , w3252 );
and ( w4134 , w4133 , w4132 );
and ( w4135 , w4134 , w6380 );
nor ( w4136 , w4135 , g3 );
and ( w4137 , w4136 , g4 );
and ( w4138 , w4137 , g10 );
and ( w4139 , w4138 , w15 );
nor ( w4140 , w4139 , w3929 );
nor ( w4141 , w4118 , w4140 );
nor ( w4142 , w4141 , g12 );
nor ( w4143 , w4142 , w3996 );
and ( w4144 , w4143 , w7097 );
and ( w4145 , w4144 , g4 );
not ( w4146 , w4145 );
and ( w4147 , w4146 , w4110 );
not ( w4148 , w4147 );
and ( w4149 , w4148 , g10 );
not ( w4150 , w4149 );
and ( w4151 , w4150 , w4064 );
nor ( w4152 , w4151 , g8 );
and ( w4153 , w4152 , w15 );
nor ( w4154 , w4153 , w3929 );
and ( w4155 , w6380 , g10 );
nor ( w4156 , w4155 , w3929 );
nor ( w4157 , w4156 , g2 );
and ( w4158 , w4157 , w7102 );
and ( w4159 , w4158 , w7183 );
and ( w4160 , w4159 , w7097 );
and ( w4161 , w4160 , w2625 );
nor ( w4162 , w4161 , w3929 );
and ( w4163 , w3668 , w7097 );
nor ( w4164 , w4163 , w3929 );
not ( w4165 , w4164 );
and ( w4166 , w4165 , g2 );
and ( w4167 , w4166 , w7102 );
not ( w4168 , w4167 );
and ( w4169 , w4168 , w4162 );
nor ( w4170 , w4169 , g10 );
not ( w4171 , w4170 );
and ( w4172 , w4171 , w4018 );
nor ( w4173 , w4172 , w15 );
and ( w4174 , w4173 , w2625 );
nor ( w4175 , w4174 , w3929 );
not ( w4176 , w3885 );
and ( w4177 , w4176 , w4175 );
nor ( w4178 , w4177 , g12 );
and ( w4179 , w4178 , w6997 );
not ( w4180 , w4179 );
and ( w4181 , w4180 , w4018 );
nor ( w4182 , w4181 , w15 );
and ( w4183 , w4182 , w7097 );
nor ( w4184 , w4183 , w3929 );
not ( w4185 , w4184 );
and ( w4186 , w4185 , w2625 );
nor ( w4187 , w4186 , w3929 );
and ( w4188 , w4162 , w4187 );
and ( w4189 , w4154 , w4188 );
and ( w4190 , w3663 , g3 );
not ( w4191 , w4190 );
and ( w4192 , w4191 , w4154 );
not ( w4193 , w4192 );
and ( w4194 , w4193 , g2 );
and ( w4195 , w15 , g3 );
nor ( w4196 , g2 , w3885 );
not ( w4197 , w4196 );
and ( w4198 , w4197 , g4 );
nor ( w4199 , w4198 , w1746 );
nor ( w4200 , g3 , w4199 );
and ( w4201 , w4200 , w6380 );
nor ( w4202 , w4201 , w3929 );
nor ( w4203 , w4202 , w15 );
and ( w4204 , w4203 , w6997 );
not ( w4205 , w4204 );
and ( w4206 , w4205 , w4054 );
not ( w4207 , w4206 );
and ( w4208 , w4207 , w8 );
not ( w4209 , w4208 );
and ( w4210 , w4154 , w4209 );
not ( w4211 , w4195 );
and ( w4212 , w4211 , w4210 );
nor ( w4213 , w4212 , g12 );
and ( w4214 , w4213 , w7213 );
and ( w4215 , w4214 , w3885 );
nor ( w4216 , w94 , g12 );
and ( w4217 , w4216 , w7183 );
and ( w4218 , w4217 , w7102 );
not ( w4219 , w4218 );
and ( w4220 , w4219 , w4154 );
not ( w4221 , w4220 );
and ( w4222 , w4221 , g10 );
nor ( w4223 , w4222 , w4208 );
not ( w4224 , w4223 );
and ( w4225 , w4224 , w8 );
nor ( w4226 , w4215 , w4225 );
not ( w4227 , w4226 );
and ( w4228 , w4227 , g10 );
nor ( w4229 , w4228 , w4208 );
not ( w4230 , w4229 );
and ( w4231 , w4230 , w8 );
nor ( w4232 , w4194 , w4231 );
not ( w4233 , w4232 );
and ( w4234 , w4233 , g4 );
nor ( w4235 , w4234 , w4225 );
not ( w4236 , w4235 );
and ( w4237 , w4236 , g10 );
nor ( w4238 , w4237 , w4208 );
not ( w4239 , w4238 );
and ( w4240 , w4239 , w8 );
not ( w4241 , w4240 );
and ( w4242 , w4189 , w4241 );
not ( w4243 , w4115 );
and ( w4244 , w4243 , w4242 );
not ( w4245 , w4244 );
and ( w4246 , w4245 , w2625 );
nor ( w4247 , w4246 , w4240 );
not ( w4248 , w4067 );
and ( w4249 , w4248 , w4247 );
not ( w4250 , w4249 );
and ( w4251 , w4250 , w2625 );
nor ( w4252 , w4251 , w4240 );
not ( w4253 , w3889 );
and ( w4254 , w4253 , w4252 );
not ( w4255 , w4254 );
and ( w4256 , w4255 , g4 );
not ( w4257 , w4256 );
and ( w4258 , w4257 , w4247 );
not ( w4259 , w4258 );
and ( w4260 , w4259 , g3 );
not ( w4261 , w4260 );
and ( w4262 , w4261 , w4242 );
not ( w4263 , w4262 );
and ( w4264 , w4263 , w2625 );
nor ( w4265 , w4264 , w4240 );
and ( t_4 , w4265 , g11 );
and ( w4266 , w7213 , g10 );
nor ( w4267 , w3885 , g10 );
nor ( w4268 , w4267 , g10 );
and ( w4269 , w4268 , w6945 );
nor ( w4270 , w3 , g6 );
and ( w4271 , w4269 , w4643 );
nor ( w4272 , w4266 , w4271 );
not ( w4273 , w4272 );
and ( w4274 , w4273 , g4 );
and ( w4275 , w148 , w4643 );
nor ( w4276 , w4266 , w4275 );
nor ( w4277 , w4276 , g4 );
and ( w4278 , w4277 , w6945 );
and ( w4279 , w4278 , w4643 );
nor ( w4280 , w4274 , w4279 );
nor ( w4281 , w4280 , g1 );
and ( w4282 , w4281 , w7183 );
and ( w4283 , w1032 , g4 );
nor ( w4284 , g2 , g1 );
and ( w4285 , w7213 , w3 );
nor ( w4286 , w3472 , g3 );
nor ( w4287 , w4285 , w4286 );
and ( w4288 , w4287 , g1 );
and ( w4289 , w4288 , g10 );
nor ( w4290 , w4289 , g3 );
and ( w4291 , w4290 , w5796 );
not ( w4292 , w4291 );
and ( w4293 , w4292 , w15 );
nor ( w4294 , w4293 , g3 );
and ( w4295 , w4344 , w4294 );
nor ( w4296 , w4295 , g4 );
and ( w4297 , w4296 , g10 );
and ( w4298 , w4297 , w4643 );
nor ( w4299 , w150 , g4 );
and ( w4300 , w4299 , g10 );
nor ( w4301 , w4300 , g3 );
and ( w4302 , w6973 , w4301 );
nor ( w4303 , w4302 , g1 );
not ( w4304 , w401 );
and ( w4305 , w4304 , g4 );
not ( w4306 , w4305 );
and ( w4307 , w4306 , g4 );
nor ( w4308 , w4294 , g4 );
not ( w4309 , w4308 );
and ( w4310 , w4309 , w4270 );
nor ( w4311 , w4310 , w3 );
nor ( w4312 , w4311 , g3 );
not ( w4313 , w4307 );
and ( w4314 , w4313 , w4312 );
not ( w4315 , w4314 );
and ( w4316 , w4315 , g1 );
and ( w4317 , w4316 , g10 );
and ( w4318 , w484 , w6945 );
and ( w4319 , w4318 , w6997 );
nor ( w4320 , g4 , w4319 );
nor ( w4321 , w4320 , g1 );
and ( w4322 , w4321 , w7183 );
and ( w4323 , w4322 , w6997 );
and ( w4324 , w4344 , g4 );
nor ( w4325 , w674 , g3 );
and ( w4326 , w4325 , w7102 );
not ( w4327 , w4326 );
and ( w4328 , w4327 , w15 );
not ( w4329 , w4324 );
and ( w4330 , w4329 , w4328 );
and ( w4331 , w4330 , w6997 );
nor ( w4332 , w4331 , g3 );
and ( w4333 , w4332 , w4933 );
and ( w4334 , w4333 , w4270 );
not ( w4335 , w4334 );
and ( w4336 , w4335 , w15 );
not ( w4337 , w4285 );
and ( w4338 , w4337 , w4336 );
and ( w4339 , w4338 , w6945 );
not ( w4340 , w4339 );
and ( w4341 , w4340 , g4 );
not ( w4342 , w4341 );
and ( w4343 , w4342 , g4 );
not ( w4344 , w4284 );
and ( w4345 , w4344 , w3 );
and ( w4346 , w4328 , w6997 );
not ( w4347 , w4345 );
and ( w4348 , w4347 , w4346 );
and ( w4349 , w4348 , w7102 );
nor ( w4350 , w4349 , g3 );
not ( w4351 , w4343 );
and ( w4352 , w4351 , w4350 );
and ( w4353 , w4352 , w6997 );
nor ( w4354 , w4353 , g10 );
nor ( w4355 , w4354 , g8 );
not ( w4356 , w4355 );
and ( w4357 , w4356 , w15 );
nor ( w4358 , w4357 , g3 );
not ( w4359 , w4323 );
and ( w4360 , w4359 , w4358 );
nor ( w4361 , w4360 , w3 );
nor ( w4362 , w4361 , g3 );
not ( w4363 , w4317 );
and ( w4364 , w4363 , w4362 );
and ( w4365 , w4364 , w4270 );
nor ( w4366 , w4365 , w3 );
nor ( w4367 , w4366 , g3 );
not ( w4368 , w4303 );
and ( w4369 , w4368 , w4367 );
not ( w4370 , w4369 );
and ( w4371 , w4370 , g10 );
not ( w4372 , w4371 );
and ( w4373 , w4372 , w4362 );
and ( w4374 , w4373 , w4933 );
and ( w4375 , w4374 , w4270 );
nor ( w4376 , w4375 , w3 );
nor ( w4377 , w4376 , g3 );
not ( w4378 , w4298 );
and ( w4379 , w4378 , w4377 );
not ( w4380 , w4283 );
and ( w4381 , w4380 , w4379 );
not ( w4382 , w4381 );
and ( w4383 , w4382 , g10 );
nor ( w4384 , w4383 , g8 );
not ( w4385 , w4384 );
and ( w4386 , w4385 , w15 );
not ( w4387 , w4386 );
and ( w4388 , w4387 , w4358 );
nor ( w4389 , w4388 , w4270 );
not ( w4390 , w4389 );
and ( w4391 , w4390 , w4377 );
not ( w4392 , w4282 );
and ( w4393 , w4392 , w4391 );
nor ( w4394 , w4393 , w4270 );
not ( w4395 , w4394 );
and ( w4396 , w4395 , w4377 );
nor ( w4397 , w4396 , g11 );
and ( w4398 , w401 , w3 );
nor ( w4399 , w4398 , w4270 );
nor ( w4400 , w3 , w4270 );
not ( w4401 , w4400 );
and ( w4402 , w4401 , g10 );
not ( w4403 , w4402 );
and ( w4404 , w4403 , g10 );
nor ( w4405 , g2 , w4404 );
nor ( w4406 , w4405 , w3 );
and ( w4407 , w4406 , g13 );
not ( w4408 , w4407 );
and ( w4409 , w4408 , g10 );
not ( w4410 , w4409 );
and ( w4411 , w4410 , g4 );
and ( w4412 , w6945 , g12 );
and ( w4413 , w4412 , w6471 );
and ( w4414 , w4413 , g10 );
not ( w4415 , w4414 );
and ( w4416 , w4415 , g11 );
and ( w4417 , w4437 , w4416 );
and ( w4418 , w4417 , w5796 );
not ( w4419 , w4418 );
and ( w4420 , w4419 , w15 );
not ( w4421 , w4420 );
and ( w4422 , w4421 , w3 );
not ( w4423 , w1906 );
and ( w4424 , w4423 , g11 );
and ( w4425 , w4424 , w7097 );
not ( w4426 , w4425 );
and ( w4427 , w4426 , g12 );
and ( w4428 , w4427 , w6945 );
not ( w4429 , w4428 );
and ( w4430 , w4429 , g10 );
not ( w4431 , w4430 );
and ( w4432 , w4431 , g10 );
and ( w4433 , w4432 , g4 );
not ( w4434 , w4433 );
and ( w4435 , w4434 , g11 );
and ( w4436 , w4435 , w7097 );
not ( w4437 , w578 );
and ( w4438 , w4437 , w4436 );
and ( w4439 , w4438 , w4270 );
not ( w4440 , w4439 );
and ( w4441 , w4440 , g2 );
and ( w4442 , w526 , w4643 );
and ( w4443 , w4442 , w6471 );
not ( w4444 , w4443 );
and ( w4445 , w4444 , g11 );
and ( w4446 , w4445 , w7097 );
not ( w4447 , w4442 );
and ( w4448 , w4447 , w4446 );
and ( w4449 , w4448 , w7213 );
nor ( w4450 , w4449 , g2 );
and ( w4451 , w4450 , w6471 );
not ( w4452 , w4451 );
and ( w4453 , w4452 , g10 );
not ( w4454 , w4453 );
and ( w4455 , w4454 , g10 );
not ( w4456 , w4455 );
and ( w4457 , w4456 , g11 );
and ( w4458 , w4457 , w7097 );
not ( w4459 , w4441 );
and ( w4460 , w4459 , w4458 );
nor ( w4461 , w4460 , g13 );
not ( w4462 , w4461 );
and ( w4463 , w4462 , g10 );
not ( w4464 , w4463 );
and ( w4465 , w4464 , g10 );
and ( w4466 , w4465 , g4 );
not ( w4467 , w4466 );
and ( w4468 , w4467 , g11 );
and ( w4469 , w4468 , w7097 );
nor ( w4470 , w4422 , w4469 );
not ( w4471 , w4470 );
and ( w4472 , w4471 , g2 );
not ( w4473 , w4472 );
and ( w4474 , w4473 , g2 );
not ( w4475 , w4474 );
and ( w4476 , w4475 , w4458 );
nor ( w4477 , w4476 , g13 );
not ( w4478 , w4477 );
and ( w4479 , w4478 , g10 );
not ( w4480 , w4479 );
and ( w4481 , w4480 , g10 );
and ( w4482 , w4481 , g4 );
not ( w4483 , w4482 );
and ( w4484 , w4483 , g11 );
and ( w4485 , w4484 , w7097 );
not ( w4486 , w4411 );
and ( w4487 , w4486 , w4485 );
not ( w4488 , w4487 );
and ( w4489 , w4488 , g10 );
nor ( w4490 , g1 , w3 );
and ( w4491 , w4490 , w6380 );
and ( w4492 , w4491 , w6997 );
not ( w4493 , w4492 );
and ( w4494 , w4493 , g11 );
not ( w4495 , w4494 );
and ( w4496 , w4495 , g13 );
not ( w4497 , w45 );
and ( w4498 , w4497 , g11 );
not ( w4499 , w4490 );
and ( w4500 , w4499 , w4498 );
nor ( w4501 , w4500 , g13 );
and ( w4502 , w4501 , w6380 );
and ( w4503 , w4502 , w6997 );
not ( w4504 , w4503 );
and ( w4505 , w4504 , g11 );
not ( w4506 , w4496 );
and ( w4507 , w4506 , w4505 );
nor ( w4508 , w4507 , w15 );
and ( w4509 , w123 , w3 );
not ( w4510 , w4509 );
and ( w4511 , w4510 , w15 );
and ( w4512 , w4511 , w4643 );
and ( w4513 , w160 , w7102 );
and ( w4514 , w4513 , w7183 );
and ( w4515 , w4284 , g4 );
nor ( w4516 , w4515 , g8 );
nor ( w4517 , w4516 , g8 );
not ( w4518 , w4517 );
and ( w4519 , w4518 , w15 );
and ( w4520 , w4519 , w6997 );
nor ( w4521 , w4520 , g10 );
not ( w4522 , w4521 );
and ( w4523 , w4522 , w4270 );
nor ( w4524 , w4523 , w3 );
not ( w4525 , w4524 );
and ( w4526 , w4525 , g11 );
and ( w4527 , w4526 , w7097 );
nor ( w4528 , w4514 , w4527 );
nor ( w4529 , w15 , w484 );
and ( w4530 , w493 , w7097 );
nor ( w4531 , w4529 , w4530 );
nor ( w4532 , w4531 , g3 );
not ( w4533 , w4532 );
and ( w4534 , w4528 , w4533 );
and ( w4535 , w4534 , w6380 );
and ( w4536 , w526 , g4 );
and ( w4537 , w6945 , w2677 );
nor ( w4538 , w150 , w3 );
and ( w4539 , w4538 , w6997 );
and ( w4540 , w484 , g10 );
nor ( w4541 , w4540 , g3 );
and ( w4542 , w4541 , w6794 );
and ( w4543 , w4542 , w5798 );
and ( w4544 , w4543 , w5796 );
and ( w4545 , w4544 , g11 );
not ( w4546 , w4545 );
and ( w4547 , w4546 , w4270 );
nor ( w4548 , w4547 , g4 );
and ( w4549 , w4548 , w6997 );
nor ( w4550 , w4549 , g8 );
nor ( w4551 , w4550 , g9 );
and ( w4552 , w4551 , w5796 );
not ( w4553 , w748 );
and ( w4554 , w4553 , w4552 );
and ( w4555 , w4554 , w6945 );
not ( w4556 , w28 );
and ( w4557 , w4556 , g2 );
not ( w4558 , w4557 );
and ( w4559 , w4558 , g2 );
and ( w4560 , w4559 , g11 );
and ( w4561 , w4560 , g12 );
and ( w4562 , w4561 , w7102 );
and ( w4563 , w4562 , w6997 );
and ( w4564 , w4563 , g1 );
nor ( w4565 , w4555 , w4564 );
nor ( w4566 , w4565 , g13 );
and ( w4567 , w4566 , g11 );
and ( w4568 , w4567 , g12 );
nor ( w4569 , w4568 , g8 );
nor ( w4570 , w4569 , g9 );
and ( w4571 , w4570 , w5796 );
nor ( w4572 , w4539 , w4571 );
and ( w4573 , w2295 , w6997 );
nor ( w4574 , w4573 , g10 );
not ( w4575 , w4572 );
and ( w4576 , w4575 , w4574 );
nor ( w4577 , w4400 , g8 );
nor ( w4578 , w4577 , g8 );
not ( w4579 , w4578 );
and ( w4580 , w4579 , g2 );
and ( w4581 , w4580 , w4270 );
and ( w4582 , w4581 , w6997 );
nor ( w4583 , w4582 , g10 );
and ( w4584 , w4576 , w4583 );
nor ( w4585 , w4537 , w4584 );
nor ( w4586 , w4585 , g4 );
and ( w4587 , w4586 , g12 );
not ( w4588 , w4587 );
and ( w4589 , w4588 , w4270 );
and ( w4590 , w4589 , g11 );
and ( w4591 , w4590 , w7097 );
not ( w4592 , w4536 );
and ( w4593 , w4592 , w4591 );
nor ( w4594 , w650 , w4571 );
nor ( w4595 , w4594 , g4 );
and ( w4596 , w4595 , w5798 );
and ( w4597 , w4596 , w5796 );
and ( w4598 , w4597 , g12 );
not ( w4599 , w4598 );
and ( w4600 , w4599 , g11 );
and ( w4601 , w4600 , w7097 );
not ( w4602 , w4515 );
and ( w4603 , w4602 , w4601 );
and ( w4604 , w4603 , w5796 );
nor ( w4605 , w4604 , g9 );
and ( w4606 , w4605 , w5796 );
and ( w4607 , w4606 , g12 );
nor ( w4608 , w4607 , g10 );
nor ( w4609 , w4608 , g10 );
not ( w4610 , w4609 );
and ( w4611 , w4610 , w4270 );
nor ( w4612 , w4611 , w3 );
not ( w4613 , w4612 );
and ( w4614 , w4613 , g11 );
and ( w4615 , w4614 , w7097 );
and ( w4616 , w4593 , w4615 );
not ( w4617 , w4616 );
and ( w4618 , w4617 , g12 );
nor ( w4619 , w4618 , g10 );
nor ( w4620 , w4619 , g10 );
not ( w4621 , w4620 );
and ( w4622 , w4621 , w4270 );
nor ( w4623 , w4622 , w3 );
not ( w4624 , w4623 );
and ( w4625 , w4624 , g11 );
and ( w4626 , w4625 , w7097 );
not ( w4627 , w4535 );
and ( w4628 , w4627 , w4626 );
not ( w4629 , w4512 );
and ( w4630 , w4629 , w4628 );
nor ( w4631 , w4630 , g12 );
not ( w4632 , w4630 );
and ( w4633 , w4632 , g12 );
and ( w4634 , w4633 , w6997 );
and ( w4635 , w4634 , g4 );
not ( w4636 , w4635 );
and ( w4637 , w4636 , g11 );
and ( w4638 , w4637 , w7097 );
not ( w4639 , w4631 );
and ( w4640 , w4639 , w4638 );
and ( w4641 , w4640 , g2 );
nor ( w4642 , w123 , w15 );
not ( w4643 , w4270 );
and ( w4644 , w4642 , w4643 );
and ( w4645 , w578 , w7183 );
not ( w4646 , w4645 );
and ( w4647 , w4646 , w4628 );
and ( w4648 , w4647 , w4270 );
nor ( w4649 , w4648 , w3 );
not ( w4650 , w4649 );
and ( w4651 , w4650 , w4628 );
nor ( w4652 , w4651 , g10 );
and ( w4653 , w4652 , g4 );
and ( w4654 , w147 , g10 );
and ( w4655 , w4654 , w7183 );
nor ( w4656 , w4655 , g4 );
not ( w4657 , w4656 );
and ( w4658 , w4657 , g11 );
and ( w4659 , w4658 , w7097 );
nor ( w4660 , g2 , w4659 );
not ( w4661 , w4660 );
and ( w4662 , w4661 , w3 );
and ( w4663 , w147 , w4270 );
and ( w4664 , w4663 , g11 );
nor ( w4665 , w160 , w4664 );
not ( w4666 , w4665 );
and ( w4667 , w4666 , w4270 );
and ( w4668 , w4667 , g10 );
nor ( w4669 , w4668 , g4 );
not ( w4670 , w4669 );
and ( w4671 , w4670 , g11 );
and ( w4672 , w4671 , w7097 );
nor ( w4673 , w4662 , w4672 );
not ( w4674 , w4673 );
and ( w4675 , w4674 , g10 );
and ( w4676 , w7213 , w4628 );
and ( w4677 , g2 , w4628 );
and ( w4678 , w4677 , w4270 );
and ( w4679 , w4678 , w6997 );
and ( w4680 , w4679 , w7183 );
nor ( w4681 , w4680 , g4 );
not ( w4682 , w4681 );
and ( w4683 , w4682 , g11 );
and ( w4684 , w4683 , w7097 );
nor ( w4685 , w4676 , w4684 );
not ( w4686 , w4685 );
and ( w4687 , w4686 , w4270 );
and ( w4688 , w4687 , w6997 );
and ( w4689 , w4688 , w7183 );
nor ( w4690 , w4285 , w4689 );
nor ( w4691 , w4690 , g1 );
nor ( w4692 , w748 , w4684 );
nor ( w4693 , w4692 , w4584 );
and ( w4694 , w4693 , g1 );
and ( w4695 , w4694 , w6997 );
and ( w4696 , w4695 , w7183 );
nor ( w4697 , w4696 , g4 );
not ( w4698 , w4697 );
and ( w4699 , w4698 , g11 );
and ( w4700 , w4699 , w7097 );
nor ( w4701 , w4691 , w4700 );
nor ( w4702 , w4701 , g10 );
nor ( w4703 , w147 , g4 );
not ( w4704 , w4703 );
and ( w4705 , w4704 , w3 );
and ( w4706 , w2137 , w6380 );
not ( w4707 , w4706 );
and ( w4708 , w4707 , w4628 );
and ( w4709 , w4708 , w4270 );
and ( w4710 , w4709 , w6997 );
and ( w4711 , w4710 , w7183 );
nor ( w4712 , w4711 , g4 );
not ( w4713 , w4712 );
and ( w4714 , w4713 , g11 );
and ( w4715 , w4714 , w7097 );
nor ( w4716 , w4705 , w4715 );
nor ( w4717 , w4716 , g10 );
and ( w4718 , w4717 , w7183 );
nor ( w4719 , w4718 , g4 );
and ( w4720 , g12 , g10 );
and ( w4721 , w4720 , w3 );
and ( w4722 , w4721 , w5796 );
nor ( w4723 , w4722 , g8 );
not ( w4724 , w4723 );
and ( w4725 , w4724 , w15 );
and ( w4726 , w4725 , g11 );
not ( w4727 , w4726 );
and ( w4728 , g1 , w4727 );
not ( w4729 , w4728 );
and ( w4730 , w4729 , g10 );
and ( w4731 , g12 , w5026 );
and ( w4732 , w4731 , w6471 );
and ( w4733 , w4732 , w6997 );
nor ( w4734 , w4733 , g8 );
not ( w4735 , w4734 );
and ( w4736 , w4735 , w15 );
and ( w4737 , w4736 , g11 );
nor ( w4738 , w4737 , g4 );
and ( w4739 , w4738 , w5796 );
not ( w4740 , w4739 );
and ( w4741 , w4740 , w15 );
and ( w4742 , w1032 , w3 );
and ( w4743 , w4742 , w5796 );
nor ( w4744 , w4743 , g8 );
not ( w4745 , w4741 );
and ( w4746 , w4745 , w4744 );
nor ( w4747 , w4746 , g10 );
nor ( w4748 , w4747 , w4726 );
and ( w4749 , w578 , w6471 );
nor ( w4750 , w4749 , w4571 );
and ( w4751 , w4750 , w4270 );
and ( w4752 , w4751 , g11 );
nor ( w4753 , w3 , w4752 );
nor ( w4754 , w4753 , g2 );
nor ( w4755 , w4754 , g4 );
not ( w4756 , w4755 );
and ( w4757 , w4756 , g11 );
nor ( w4758 , w4678 , w4757 );
nor ( w4759 , w4758 , w4584 );
and ( w4760 , w4759 , g1 );
not ( w4761 , w4760 );
and ( w4762 , w4761 , w4744 );
nor ( w4763 , w4762 , g10 );
nor ( w4764 , w4763 , g4 );
and ( w4765 , w4764 , w5796 );
not ( w4766 , w4765 );
and ( w4767 , w4766 , w15 );
and ( w4768 , w4767 , g11 );
and ( w4769 , w4768 , w7097 );
not ( w4770 , w4769 );
and ( w4771 , w4748 , w4770 );
not ( w4772 , w4771 );
and ( w4773 , w4772 , g2 );
and ( w4774 , g1 , g10 );
nor ( w4775 , w4737 , w4769 );
and ( w4776 , w4775 , g2 );
not ( w4777 , w650 );
and ( w4778 , w4750 , w4777 );
and ( w4779 , w4778 , w6997 );
nor ( w4780 , w242 , w4779 );
nor ( w4781 , w4780 , g2 );
nor ( w4782 , w4781 , g2 );
and ( w4783 , w4782 , w4544 );
not ( w4784 , w4783 );
and ( w4785 , w4784 , g11 );
and ( w4786 , w4785 , w7097 );
not ( w4787 , w4776 );
and ( w4788 , w4787 , w4786 );
not ( w4789 , w4788 );
and ( w4790 , w4789 , w4544 );
not ( w4791 , w4790 );
and ( w4792 , w4791 , w4270 );
nor ( w4793 , w4792 , g4 );
nor ( w4794 , w4793 , g8 );
nor ( w4795 , w4794 , g8 );
not ( w4796 , w4795 );
and ( w4797 , w4796 , w15 );
and ( w4798 , w4797 , g11 );
and ( w4799 , w4798 , w7097 );
not ( w4800 , w4799 );
and ( w4801 , w4775 , w4800 );
and ( w4802 , w4801 , w7102 );
and ( w4803 , w4802 , w5796 );
not ( w4804 , w4803 );
and ( w4805 , w4804 , w15 );
nor ( w4806 , w4774 , w4805 );
nor ( w4807 , w4806 , g2 );
and ( w4808 , w4807 , w3 );
nor ( w4809 , w4808 , w4799 );
and ( w4810 , w4809 , w7102 );
nor ( w4811 , w4810 , g8 );
nor ( w4812 , w4811 , g8 );
not ( w4813 , w4812 );
and ( w4814 , w4813 , w15 );
and ( w4815 , w4814 , g11 );
and ( w4816 , w4815 , w7097 );
nor ( w4817 , w4773 , w4816 );
not ( w4818 , w4817 );
and ( w4819 , w4818 , w3 );
nor ( w4820 , w4819 , w4799 );
and ( w4821 , w4820 , w7102 );
nor ( w4822 , w4821 , g8 );
nor ( w4823 , w4822 , g8 );
not ( w4824 , w4823 );
and ( w4825 , w4824 , w15 );
and ( w4826 , w4825 , g11 );
and ( w4827 , w4826 , w7097 );
nor ( w4828 , w4730 , w4827 );
not ( w4829 , w4828 );
and ( w4830 , w4829 , g2 );
nor ( w4831 , w4830 , w4816 );
not ( w4832 , w4831 );
and ( w4833 , w4832 , w3 );
nor ( w4834 , w4833 , w4799 );
and ( w4835 , w4834 , w7102 );
nor ( w4836 , w4835 , g8 );
nor ( w4837 , w4836 , g8 );
not ( w4838 , w4837 );
and ( w4839 , w4838 , w15 );
and ( w4840 , w4839 , g11 );
and ( w4841 , w4840 , w7097 );
and ( w4842 , w4719 , w4856 );
not ( w4843 , w4842 );
and ( w4844 , w4843 , g11 );
and ( w4845 , w4844 , w7097 );
nor ( w4846 , w4702 , w4845 );
nor ( w4847 , w4846 , w15 );
nor ( w4848 , w4847 , g4 );
and ( w4849 , w4848 , w4856 );
not ( w4850 , w4849 );
and ( w4851 , w4850 , g11 );
and ( w4852 , w4851 , w7097 );
nor ( w4853 , w4675 , w4852 );
nor ( w4854 , w4853 , w15 );
nor ( w4855 , w4854 , g4 );
not ( w4856 , w4841 );
and ( w4857 , w4855 , w4856 );
not ( w4858 , w4857 );
and ( w4859 , w4858 , g11 );
and ( w4860 , w4859 , w7097 );
not ( w4861 , w4653 );
and ( w4862 , w4861 , w4860 );
not ( w4863 , w4644 );
and ( w4864 , w4863 , w4862 );
and ( w4865 , w4864 , w7213 );
nor ( w4866 , w4865 , g10 );
and ( w4867 , w4866 , g4 );
not ( w4868 , w4867 );
and ( w4869 , w4868 , w4860 );
nor ( w4870 , w4641 , w4869 );
and ( w4871 , w4870 , w6997 );
and ( w4872 , w4871 , g4 );
not ( w4873 , w4872 );
and ( w4874 , w4873 , w4860 );
not ( w4875 , w4508 );
and ( w4876 , w4875 , w4874 );
and ( w4877 , w4876 , w4638 );
and ( w4878 , w4877 , g2 );
nor ( w4879 , w4878 , w4869 );
nor ( w4880 , w4489 , w4879 );
not ( w4881 , w4399 );
and ( w4882 , w4881 , w4880 );
nor ( w4883 , w4882 , g1 );
not ( w4884 , w4883 );
and ( w4885 , w4884 , g10 );
not ( w4886 , w4885 );
and ( w4887 , w4886 , g4 );
not ( w4888 , w4887 );
and ( w4889 , w4888 , w4485 );
not ( w4890 , w4889 );
and ( w4891 , w4890 , g10 );
nor ( w4892 , w4891 , w4879 );
nor ( w4893 , w2677 , w4892 );
and ( w4894 , w4893 , w6535 );
not ( w4895 , w4894 );
and ( w4896 , w4895 , w3 );
nor ( w4897 , w4896 , w4270 );
not ( w4898 , w4897 );
and ( w4899 , w4898 , w4880 );
nor ( w4900 , w4899 , g1 );
and ( w4901 , w4900 , g13 );
not ( w4902 , w4901 );
and ( w4903 , w4902 , g10 );
not ( w4904 , w4903 );
and ( w4905 , w4904 , g4 );
not ( w4906 , w4905 );
and ( w4907 , w4906 , w4485 );
not ( w4908 , w4907 );
and ( w4909 , w4908 , g10 );
nor ( w4910 , w4909 , w4879 );
not ( w4911 , w4910 );
and ( w4912 , w4911 , g11 );
nor ( w4913 , w4912 , g3 );
not ( w4914 , w4397 );
and ( w4915 , w4914 , w4913 );
nor ( w4916 , g3 , w4915 );
nor ( w4917 , g1 , w4915 );
nor ( w4918 , w4917 , w4916 );
and ( w4919 , w4918 , w7213 );
not ( w4920 , w4919 );
and ( w4921 , w4920 , g4 );
nor ( w4922 , w4921 , w4916 );
nor ( w4923 , w1032 , w4922 );
and ( w4924 , w4923 , w5698 );
nor ( w4925 , w4924 , w4916 );
nor ( w4926 , w4925 , w15 );
and ( w4927 , w5668 , g2 );
and ( w4928 , w4918 , g10 );
and ( w4929 , g1 , w5698 );
and ( w4930 , w4929 , g4 );
nor ( w4931 , w4930 , w4916 );
and ( w4932 , w4931 , w6997 );
not ( w4933 , g6 );
and ( w4934 , w4932 , w4933 );
and ( w4935 , w4934 , w4270 );
nor ( w4936 , w4935 , w4915 );
and ( w4937 , w5438 , w4936 );
and ( w4938 , w4937 , w7094 );
nor ( w4939 , w4938 , w4916 );
and ( w4940 , w4939 , w4270 );
nor ( w4941 , w4940 , w4915 );
nor ( w4942 , w4941 , g2 );
nor ( w4943 , w4942 , g2 );
nor ( w4944 , w4943 , w4916 );
nor ( w4945 , w4918 , g4 );
nor ( w4946 , w4945 , w4916 );
nor ( w4947 , w4946 , w15 );
nor ( w4948 , w4947 , w4916 );
and ( w4949 , w5668 , g1 );
nor ( w4950 , w4949 , w4270 );
nor ( w4951 , w4950 , w4916 );
nor ( w4952 , w4951 , w4915 );
not ( w4953 , w4952 );
and ( w4954 , w4953 , g2 );
not ( w4955 , w4954 );
and ( w4956 , w4955 , g2 );
and ( w4957 , w5668 , w3 );
and ( w4958 , w4918 , w4270 );
nor ( w4959 , w4958 , w4915 );
and ( w4960 , w4959 , w7183 );
not ( w4961 , w4957 );
and ( w4962 , w4961 , w4960 );
nor ( w4963 , w4962 , w4916 );
nor ( w4964 , w4963 , g2 );
nor ( w4965 , w4964 , w4916 );
not ( w4966 , w4965 );
and ( w4967 , w4966 , g4 );
nor ( w4968 , w4967 , w4916 );
not ( w4969 , w4956 );
and ( w4970 , w4969 , w4968 );
not ( w4971 , w4970 );
and ( w4972 , w4971 , g4 );
and ( w4973 , w4918 , g2 );
nor ( w4974 , w4919 , w4915 );
and ( w4975 , w4974 , w7102 );
nor ( w4976 , w4975 , w4916 );
not ( w4977 , w4976 );
and ( w4978 , w4977 , g10 );
nor ( w4979 , w4978 , w4916 );
nor ( w4980 , w4979 , w15 );
nor ( w4981 , w4980 , w4916 );
nor ( w4982 , w4973 , w4981 );
and ( w4983 , w4982 , w6535 );
nor ( w4984 , w4983 , w4916 );
and ( w4985 , w4984 , w3 );
nor ( w4986 , w4985 , w4270 );
and ( w4987 , w5346 , g2 );
nor ( w4988 , w4987 , w4916 );
and ( w4989 , w4988 , w4270 );
nor ( w4990 , w4989 , w3 );
nor ( w4991 , w4990 , w4916 );
nor ( w4992 , w4991 , g4 );
nor ( w4993 , w4992 , w4916 );
nor ( w4994 , w4993 , w15 );
nor ( w4995 , w4994 , w4916 );
not ( w4996 , w4986 );
and ( w4997 , w4996 , w4995 );
not ( w4998 , w4997 );
and ( w4999 , w4998 , g10 );
nor ( w5000 , w4999 , w4916 );
not ( w5001 , w5000 );
and ( w5002 , w5001 , g12 );
nor ( w5003 , w4972 , w5002 );
and ( w5004 , w5003 , w5668 );
not ( w5005 , w5004 );
and ( w5006 , w5005 , g10 );
nor ( w5007 , w5006 , w4916 );
nor ( w5008 , w4957 , w4270 );
nor ( w5009 , w5008 , g10 );
nor ( w5010 , w4918 , w15 );
nor ( w5011 , w4916 , g8 );
nor ( w5012 , w5011 , g8 );
nor ( w5013 , w5010 , w5012 );
not ( w5014 , w5013 );
and ( w5015 , w5014 , g13 );
nor ( w5016 , w4918 , g13 );
nor ( w5017 , w5016 , w4916 );
nor ( w5018 , w5017 , w15 );
nor ( w5019 , w5018 , w4916 );
and ( w5020 , w4988 , w3 );
nor ( w5021 , w5020 , w4270 );
nor ( w5022 , w5021 , w4916 );
not ( w5023 , w5022 );
and ( w5024 , w5023 , g4 );
nor ( w5025 , w5024 , w4916 );
not ( w5026 , w4571 );
and ( w5027 , w5025 , w5026 );
and ( w5028 , w5027 , w6997 );
nor ( w5029 , w5028 , g10 );
and ( w5030 , w5029 , w6471 );
and ( w5031 , w5030 , g12 );
nor ( w5032 , w5031 , w4916 );
and ( w5033 , w5032 , w5796 );
not ( w5034 , w5033 );
and ( w5035 , w5034 , w15 );
nor ( w5036 , w5035 , w4916 );
and ( w5037 , w5019 , w5036 );
nor ( w5038 , w5037 , w3 );
and ( w5039 , w5038 , g12 );
nor ( w5040 , w5039 , w4916 );
not ( w5041 , w5040 );
and ( w5042 , w5041 , g4 );
not ( w5043 , w4949 );
and ( w5044 , w5043 , g13 );
and ( w5045 , w6127 , g11 );
nor ( w5046 , g12 , w5045 );
and ( w5047 , w4917 , g12 );
nor ( w5048 , w5046 , w5047 );
nor ( w5049 , w5048 , w4915 );
and ( w5050 , w5049 , w6471 );
nor ( w5051 , w5050 , w4916 );
not ( w5052 , w5044 );
and ( w5053 , w5052 , w5051 );
nor ( w5054 , w5053 , w4915 );
and ( w5055 , w5054 , g4 );
nor ( w5056 , w5055 , w4916 );
nor ( w5057 , w5056 , w15 );
nor ( w5058 , w5057 , w4916 );
and ( w5059 , w4918 , w6997 );
nor ( w5060 , w5059 , w4915 );
and ( w5061 , w5060 , w7213 );
not ( w5062 , w5061 );
and ( w5063 , w5062 , w3 );
nor ( w5064 , w5063 , w4915 );
nor ( w5065 , w5064 , w4916 );
nor ( w5066 , w5065 , g4 );
nor ( w5067 , w5066 , w4916 );
and ( w5068 , w5067 , w3 );
nor ( w5069 , w5068 , w4915 );
and ( w5070 , w5069 , w7213 );
nor ( w5071 , w5070 , w4916 );
and ( w5072 , w5071 , w6997 );
and ( w5073 , w5072 , w5796 );
not ( w5074 , w5073 );
and ( w5075 , w5074 , w15 );
nor ( w5076 , w5075 , w4916 );
and ( w5077 , w5076 , w3 );
and ( w5078 , w5077 , w6997 );
and ( w5079 , w5058 , w5078 );
nor ( w5080 , w5079 , w4915 );
and ( w5081 , w5080 , w6535 );
not ( w5082 , w5081 );
and ( w5083 , w5082 , w3 );
nor ( w5084 , w4931 , w3 );
nor ( w5085 , w5084 , w4916 );
nor ( w5086 , w5085 , g10 );
nor ( w5087 , w5086 , w4916 );
and ( w5088 , w5087 , w7213 );
nor ( w5089 , w5088 , g2 );
nor ( w5090 , w5089 , w4916 );
not ( w5091 , w5090 );
and ( w5092 , w5091 , g12 );
nor ( w5093 , w5092 , w4916 );
not ( w5094 , w5093 );
and ( w5095 , w5094 , g13 );
and ( w5096 , w78 , w6471 );
not ( w5097 , w5096 );
and ( w5098 , w5097 , w5036 );
not ( w5099 , w5098 );
and ( w5100 , w5099 , g11 );
nor ( w5101 , w5095 , w5100 );
nor ( w5102 , w5101 , w4915 );
nor ( w5103 , w5102 , w4916 );
not ( w5104 , w5103 );
and ( w5105 , w15 , w5104 );
nor ( w5106 , w5105 , w4916 );
not ( w5107 , w5106 );
and ( w5108 , w5107 , g4 );
nor ( w5109 , w5108 , w4916 );
nor ( w5110 , w4949 , w15 );
and ( w5111 , w5110 , w6997 );
and ( w5112 , w5111 , w6794 );
and ( w5113 , w5112 , w5698 );
and ( w5114 , w5113 , w7102 );
nor ( w5115 , w5114 , w4916 );
and ( w5116 , w5115 , w7213 );
nor ( w5117 , w5116 , g2 );
nor ( w5118 , w5117 , w4916 );
and ( w5119 , w5698 , g2 );
and ( w5120 , w5119 , w15 );
and ( w5121 , w484 , g3 );
not ( w5122 , w5121 );
and ( w5123 , w5122 , g3 );
nor ( w5124 , w5123 , w4544 );
and ( w5125 , w5124 , w5796 );
nor ( w5126 , w5125 , g8 );
and ( w5127 , w5120 , w5126 );
not ( w5128 , w5127 );
and ( w5129 , w5118 , w5128 );
and ( w5130 , w5129 , w6997 );
nor ( w5131 , w5130 , g10 );
not ( w5132 , w5131 );
and ( w5133 , w5132 , w4270 );
nor ( w5134 , w5133 , w3 );
and ( w5135 , w5134 , w7102 );
not ( w5136 , w5135 );
and ( w5137 , w5109 , w5136 );
and ( w5138 , w5137 , w4270 );
nor ( w5139 , w5138 , w4915 );
nor ( w5140 , w5139 , g2 );
nor ( w5141 , w5140 , g2 );
nor ( w5142 , w5141 , w4916 );
and ( w5143 , w5142 , w6997 );
nor ( w5144 , w5143 , g10 );
and ( w5145 , w5144 , g11 );
not ( w5146 , w5083 );
and ( w5147 , w5146 , w5145 );
nor ( w5148 , w5147 , w4916 );
not ( w5149 , w5042 );
and ( w5150 , w5149 , w5148 );
and ( w5151 , w5150 , g2 );
not ( w5152 , w5151 );
and ( w5153 , w5152 , g2 );
nor ( w5154 , w5153 , w5147 );
and ( w5155 , w5154 , w5668 );
nor ( w5156 , w5155 , g10 );
nor ( w5157 , w5156 , w4916 );
not ( w5158 , w5157 );
and ( w5159 , w5158 , g11 );
nor ( w5160 , w5015 , w5159 );
and ( w5161 , w5160 , w5668 );
and ( w5162 , w5161 , w4270 );
nor ( w5163 , w5162 , w3 );
nor ( w5164 , w5163 , w4916 );
not ( w5165 , w5164 );
and ( w5166 , w5165 , g4 );
nor ( w5167 , w5166 , w4916 );
and ( w5168 , w5167 , w5148 );
and ( w5169 , w5168 , g2 );
not ( w5170 , w5169 );
and ( w5171 , w5170 , g2 );
nor ( w5172 , w5171 , w5147 );
and ( w5173 , w5172 , w5668 );
and ( w5174 , w5173 , w6997 );
nor ( w5175 , w5174 , g10 );
and ( w5176 , w5175 , g11 );
not ( w5177 , w5176 );
and ( w5178 , w5009 , w5177 );
and ( w5179 , w5178 , w5148 );
nor ( w5180 , w5179 , g10 );
nor ( w5181 , w5180 , w4916 );
not ( w5182 , w4412 );
and ( w5183 , w5182 , g11 );
and ( w5184 , w5183 , w5668 );
and ( w5185 , w5184 , w7213 );
nor ( w5186 , w5185 , g2 );
and ( w5187 , w5186 , w5698 );
nor ( w5188 , w5187 , w4916 );
not ( w5189 , w5188 );
and ( w5190 , w5189 , g10 );
nor ( w5191 , w4987 , g10 );
and ( w5192 , w5191 , w5616 );
nor ( w5193 , w5192 , g10 );
nor ( w5194 , w5193 , w4916 );
and ( w5195 , w5194 , w3 );
nor ( w5196 , w5195 , w4915 );
and ( w5197 , w5196 , g4 );
nor ( w5198 , w5197 , w4916 );
not ( w5199 , w5198 );
and ( w5200 , w5199 , g12 );
and ( w5201 , w5200 , g11 );
nor ( w5202 , w5190 , w5201 );
and ( w5203 , w5202 , w5668 );
and ( w5204 , w5203 , w3 );
nor ( w5205 , w5204 , w4270 );
nor ( w5206 , w4918 , g2 );
nor ( w5207 , w5206 , w4916 );
and ( w5208 , w5207 , w4270 );
not ( w5209 , w5208 );
and ( w5210 , w5209 , g10 );
and ( w5211 , w5210 , w6794 );
nor ( w5212 , w5211 , w5176 );
and ( w5213 , w5212 , w5668 );
not ( w5214 , w5213 );
and ( w5215 , w5214 , g4 );
and ( w5216 , w5215 , g13 );
nor ( w5217 , w5216 , w4916 );
not ( w5218 , w5217 );
and ( w5219 , w5218 , g12 );
and ( w5220 , w5219 , g11 );
nor ( w5221 , w5205 , w5220 );
and ( w5222 , w5221 , w5668 );
not ( w5223 , w5222 );
and ( w5224 , w5223 , g4 );
and ( w5225 , w4973 , w3 );
not ( w5226 , w5225 );
and ( w5227 , w5226 , g2 );
nor ( w5228 , w5227 , w4916 );
not ( w5229 , w5228 );
and ( w5230 , w5229 , g10 );
nor ( w5231 , w5230 , g4 );
nor ( w5232 , w5231 , w4270 );
and ( w5233 , w5232 , w7102 );
and ( w5234 , w5668 , g10 );
not ( w5235 , w5234 );
and ( w5236 , w5235 , w5066 );
nor ( w5237 , w5236 , w4916 );
nor ( w5238 , w5237 , g2 );
nor ( w5239 , w5238 , w4916 );
nor ( w5240 , w5239 , w4270 );
nor ( w5241 , w5240 , w4916 );
and ( w5242 , w5241 , w5796 );
not ( w5243 , w5242 );
and ( w5244 , w5243 , w15 );
nor ( w5245 , w5244 , w4916 );
not ( w5246 , w5233 );
and ( w5247 , w5246 , w5245 );
and ( w5248 , w5300 , g2 );
nor ( w5249 , w4916 , g10 );
nor ( w5250 , w5249 , g10 );
and ( w5251 , w4945 , w6794 );
and ( w5252 , w5251 , g10 );
nor ( w5253 , w5250 , w5252 );
and ( w5254 , w5253 , w5668 );
and ( w5255 , w5254 , w7213 );
nor ( w5256 , w5255 , g2 );
nor ( w5257 , w5256 , w4916 );
not ( w5258 , w5257 );
and ( w5259 , w5258 , w15 );
nor ( w5260 , w5248 , w5259 );
and ( w5261 , w5260 , w5668 );
and ( w5262 , w5261 , w5093 );
not ( w5263 , w5262 );
and ( w5264 , w5263 , g13 );
nor ( w5265 , w5264 , w4916 );
and ( w5266 , w5265 , w5796 );
not ( w5267 , w5266 );
and ( w5268 , w5267 , w15 );
nor ( w5269 , w5268 , w4916 );
and ( w5270 , w5247 , w5269 );
and ( w5271 , w5270 , w5148 );
and ( w5272 , w5271 , w5093 );
not ( w5273 , w5272 );
and ( w5274 , w5273 , g13 );
nor ( w5275 , w5274 , w4916 );
and ( w5276 , w5275 , w5796 );
not ( w5277 , w5276 );
and ( w5278 , w5277 , w15 );
nor ( w5279 , w4988 , g4 );
nor ( w5280 , w5279 , w4916 );
and ( w5281 , w5187 , g4 );
nor ( w5282 , w5281 , w4916 );
not ( w5283 , w5282 );
and ( w5284 , w5283 , g10 );
nor ( w5285 , w5284 , w4916 );
and ( w5286 , w5280 , w5285 );
and ( w5287 , w5286 , w3 );
nor ( w5288 , w5287 , w4270 );
and ( w5289 , w5346 , g4 );
nor ( w5290 , w5289 , w5252 );
and ( w5291 , w5290 , w7213 );
and ( w5292 , w5291 , w5668 );
nor ( w5293 , w5292 , w4915 );
and ( w5294 , w5293 , w6794 );
nor ( w5295 , w5294 , w4916 );
not ( w5296 , w5295 );
and ( w5297 , w5296 , g10 );
and ( w5298 , w5297 , w6471 );
and ( w5299 , w5298 , g12 );
not ( w5300 , w4927 );
and ( w5301 , w5300 , w5299 );
nor ( w5302 , w5301 , w4916 );
not ( w5303 , w5288 );
and ( w5304 , w5303 , w5302 );
not ( w5305 , w5304 );
and ( w5306 , w5305 , g10 );
nor ( w5307 , w5306 , w4916 );
and ( w5308 , w5307 , w5036 );
nor ( w5309 , w5308 , g13 );
and ( w5310 , w5309 , g12 );
nor ( w5311 , w5310 , w4916 );
and ( w5312 , w5311 , w5796 );
not ( w5313 , w5312 );
and ( w5314 , w5313 , w15 );
nor ( w5315 , w5314 , w4916 );
not ( w5316 , w5278 );
and ( w5317 , w5316 , w5315 );
not ( w5318 , w5317 );
and ( w5319 , w5318 , g12 );
and ( w5320 , w5319 , g11 );
nor ( w5321 , w5224 , w5320 );
and ( w5322 , w5321 , w5093 );
not ( w5323 , w5322 );
and ( w5324 , w5323 , g13 );
nor ( w5325 , w5324 , w4916 );
and ( w5326 , w5325 , w5796 );
not ( w5327 , w5326 );
and ( w5328 , w5327 , w15 );
nor ( w5329 , w5328 , w4916 );
and ( w5330 , w5329 , w5315 );
not ( w5331 , w5330 );
and ( w5332 , w5331 , g11 );
and ( w5333 , w5181 , w5337 );
and ( w5334 , w5007 , w5333 );
nor ( w5335 , w5334 , w15 );
nor ( w5336 , w5335 , w4916 );
not ( w5337 , w5332 );
and ( w5338 , w5336 , w5337 );
not ( w5339 , w5338 );
and ( w5340 , w5339 , g11 );
nor ( w5341 , w4916 , w5340 );
and ( w5342 , w4948 , w5341 );
and ( w5343 , w5342 , g2 );
not ( w5344 , w5343 );
and ( w5345 , w5344 , g2 );
not ( w5346 , w4918 );
and ( w5347 , w5346 , w15 );
nor ( w5348 , w5347 , w4916 );
nor ( w5349 , w5348 , g12 );
nor ( w5350 , w5349 , w5340 );
not ( w5351 , w5350 );
and ( w5352 , w5351 , g11 );
nor ( w5353 , w5010 , w5352 );
and ( w5354 , w5353 , w5668 );
not ( w5355 , w5354 );
and ( w5356 , w5355 , g4 );
and ( w5357 , w4963 , g2 );
not ( w5358 , w5357 );
and ( w5359 , w5358 , g2 );
nor ( w5360 , w5359 , g10 );
and ( w5361 , w5360 , w5668 );
nor ( w5362 , w5361 , g10 );
and ( w5363 , w5362 , w6380 );
nor ( w5364 , w5363 , w4916 );
not ( w5365 , w5364 );
and ( w5366 , w5365 , g4 );
nor ( w5367 , w5366 , w4916 );
and ( w5368 , w5367 , g2 );
not ( w5369 , w5368 );
and ( w5370 , w5369 , g2 );
nor ( w5371 , w5370 , g10 );
and ( w5372 , w5371 , w5148 );
nor ( w5373 , w5372 , g10 );
nor ( w5374 , w5373 , w5340 );
not ( w5375 , w5374 );
and ( w5376 , w5375 , g11 );
nor ( w5377 , w5376 , w4916 );
and ( w5378 , w5261 , w5377 );
not ( w5379 , w5378 );
and ( w5380 , w5379 , g11 );
nor ( w5381 , w5380 , w4916 );
not ( w5382 , w5356 );
and ( w5383 , w5382 , w5381 );
nor ( w5384 , w5383 , g2 );
nor ( w5385 , w5384 , w4916 );
not ( w5386 , w5385 );
and ( w5387 , w5386 , g10 );
not ( w5388 , w5387 );
and ( w5389 , w5388 , w5377 );
nor ( w5390 , w5389 , g12 );
nor ( w5391 , w5390 , w5340 );
not ( w5392 , w5391 );
and ( w5393 , w5392 , g11 );
nor ( w5394 , w5393 , w4916 );
and ( w5395 , w5394 , w4270 );
not ( w5396 , w5345 );
and ( w5397 , w5396 , w5395 );
nor ( w5398 , w5397 , w4915 );
and ( w5399 , w5398 , g10 );
not ( w5400 , w5399 );
and ( w5401 , w5400 , w5377 );
nor ( w5402 , w5401 , g12 );
nor ( w5403 , w5402 , w5340 );
not ( w5404 , w5403 );
and ( w5405 , w5404 , g11 );
nor ( w5406 , w5405 , w4916 );
and ( w5407 , w5406 , w4270 );
and ( w5408 , w4944 , w5407 );
nor ( w5409 , w5408 , w4915 );
nor ( w5410 , w5409 , g2 );
nor ( w5411 , w5410 , w4915 );
and ( w5412 , w5411 , w15 );
nor ( w5413 , w5412 , w4916 );
and ( w5414 , w5413 , g10 );
not ( w5415 , w5414 );
and ( w5416 , w5415 , g10 );
nor ( w5417 , w240 , w4916 );
nor ( w5418 , w5417 , w4915 );
nor ( w5419 , w5418 , g2 );
nor ( w5420 , w5419 , g10 );
not ( w5421 , w4973 );
and ( w5422 , w5421 , w5420 );
nor ( w5423 , w5422 , w4916 );
nor ( w5424 , w5423 , w15 );
nor ( w5425 , g1 , w4916 );
nor ( w5426 , w5425 , w4915 );
not ( w5427 , w5426 );
and ( w5428 , w5427 , g2 );
not ( w5429 , w5428 );
and ( w5430 , w5429 , g2 );
not ( w5431 , w5430 );
and ( w5432 , w5431 , w5408 );
nor ( w5433 , w5432 , w4915 );
and ( w5434 , w5433 , w15 );
nor ( w5435 , w5434 , w4916 );
not ( w5436 , w5435 );
and ( w5437 , w5436 , g4 );
not ( w5438 , w4928 );
and ( w5439 , w5438 , g10 );
nor ( w5440 , w5439 , w240 );
and ( w5441 , w5440 , w5668 );
nor ( w5442 , w5441 , w4915 );
not ( w5443 , w5442 );
and ( w5444 , w5443 , g2 );
not ( w5445 , w5444 );
and ( w5446 , w5445 , g2 );
nor ( w5447 , w4949 , g10 );
nor ( w5448 , w5447 , w4916 );
nor ( w5449 , w5448 , w4915 );
nor ( w5450 , w5449 , g2 );
nor ( w5451 , w5450 , g2 );
nor ( w5452 , w5451 , w4916 );
and ( w5453 , w5452 , w7102 );
nor ( w5454 , w5453 , g4 );
nor ( w5455 , w5454 , w4916 );
not ( w5456 , w5446 );
and ( w5457 , w5456 , w5455 );
nor ( w5458 , w5457 , w15 );
not ( w5459 , w5433 );
and ( w5460 , w5459 , g10 );
not ( w5461 , w5460 );
and ( w5462 , w5461 , g10 );
nor ( w5463 , w5462 , w4916 );
and ( w5464 , w5463 , w5796 );
not ( w5465 , w5464 );
and ( w5466 , w5465 , w15 );
nor ( w5467 , w5466 , w4916 );
and ( w5468 , w5467 , w7102 );
nor ( w5469 , w5468 , g4 );
and ( w5470 , w5469 , w7094 );
not ( w5471 , w5470 );
and ( w5472 , w5471 , w5407 );
not ( w5473 , w5458 );
and ( w5474 , w5473 , w5472 );
nor ( w5475 , w5474 , w4915 );
nor ( w5476 , w5475 , g4 );
nor ( w5477 , w5476 , g4 );
and ( w5478 , w5477 , w7094 );
not ( w5479 , w5478 );
and ( w5480 , w5479 , w5407 );
not ( w5481 , w5437 );
and ( w5482 , w5481 , w5480 );
nor ( w5483 , w5482 , g11 );
not ( w5484 , w5483 );
and ( w5485 , w5484 , w5407 );
not ( w5486 , w5424 );
and ( w5487 , w5486 , w5485 );
nor ( w5488 , w5487 , w4915 );
and ( w5489 , w5488 , w6997 );
nor ( w5490 , w5489 , w4916 );
not ( w5491 , w5490 );
and ( w5492 , w5491 , g4 );
not ( w5493 , w5492 );
and ( w5494 , w5493 , w5480 );
nor ( w5495 , w5494 , g11 );
not ( w5496 , w5495 );
and ( w5497 , w5496 , w5407 );
not ( w5498 , w5416 );
and ( w5499 , w5498 , w5497 );
nor ( w5500 , w5499 , w4915 );
and ( w5501 , w5500 , g4 );
not ( w5502 , w5501 );
and ( w5503 , w5502 , w5480 );
nor ( w5504 , w4927 , w5503 );
not ( w5505 , w5504 );
and ( w5506 , w5505 , w5497 );
not ( w5507 , w4926 );
and ( w5508 , w5507 , w5506 );
nor ( w5509 , w5508 , w4915 );
not ( w5510 , w5509 );
and ( w5511 , w5510 , g10 );
not ( w5512 , w5511 );
and ( w5513 , w5512 , g10 );
not ( w5514 , w5513 );
and ( w5515 , w5514 , w5497 );
nor ( w5516 , w5515 , g11 );
not ( w5517 , w5516 );
and ( w5518 , w5517 , w5407 );
nor ( w5519 , w3 , w5518 );
nor ( w5520 , w4916 , w5519 );
and ( w5521 , w5520 , g10 );
nor ( w5522 , w5518 , w4915 );
not ( w5523 , w5521 );
and ( w5524 , w5523 , w5522 );
and ( w5525 , w5524 , w6945 );
not ( w5526 , w5525 );
and ( w5527 , w5526 , w5520 );
and ( w5528 , w5527 , g4 );
and ( w5529 , w5522 , g10 );
not ( w5530 , w5529 );
and ( w5531 , w5530 , w5520 );
nor ( w5532 , w5531 , g1 );
and ( w5533 , w5524 , g1 );
not ( w5534 , w5533 );
and ( w5535 , w5534 , w5520 );
nor ( w5536 , w5535 , g11 );
nor ( w5537 , w5536 , w4916 );
not ( w5538 , w5532 );
and ( w5539 , w5538 , w5537 );
and ( w5540 , w5539 , w5520 );
and ( w5541 , w5540 , w7102 );
nor ( w5542 , w5541 , g11 );
not ( w5543 , w5542 );
and ( w5544 , w5543 , w5520 );
nor ( w5545 , w5544 , w5518 );
and ( w5546 , w5545 , w5522 );
not ( w5547 , w5528 );
and ( w5548 , w5547 , w5546 );
and ( w5549 , w5548 , w7094 );
and ( w5550 , w4917 , w5522 );
and ( w5551 , w5520 , w5148 );
and ( w5552 , w5551 , w5572 );
not ( w5553 , w5550 );
and ( w5554 , w5553 , w5552 );
nor ( w5555 , w5554 , g10 );
nor ( w5556 , w5555 , w5519 );
not ( w5557 , w5556 );
and ( w5558 , w5557 , g4 );
and ( w5559 , w5584 , g10 );
and ( w5560 , w5559 , w7102 );
nor ( w5561 , w5560 , w5519 );
and ( w5562 , w5561 , w5148 );
nor ( w5563 , w5562 , g12 );
nor ( w5564 , w5563 , w5519 );
and ( w5565 , w5564 , w5668 );
and ( w5566 , w5565 , w5572 );
not ( w5567 , w5558 );
and ( w5568 , w5567 , w5566 );
nor ( w5569 , w5568 , g12 );
not ( w5570 , w5569 );
and ( w5571 , w5570 , w5520 );
not ( w5572 , w5340 );
and ( w5573 , w5571 , w5572 );
not ( w5574 , w5573 );
and ( w5575 , w5574 , g11 );
nor ( w5576 , w5575 , w4916 );
and ( w5577 , w5576 , w5744 );
not ( w5578 , w5577 );
and ( w5579 , w5578 , w15 );
nor ( w5580 , w5549 , w5579 );
and ( w5581 , w5580 , w5744 );
and ( w5582 , w5581 , w5520 );
and ( w5583 , w5582 , g2 );
not ( w5584 , w5554 );
and ( w5585 , w5584 , g4 );
nor ( w5586 , w5585 , w4916 );
nor ( w5587 , w5586 , g11 );
and ( w5588 , w5522 , g4 );
not ( w5589 , w5588 );
and ( w5590 , w5589 , w5520 );
nor ( w5591 , w5590 , g1 );
not ( w5592 , w5591 );
and ( w5593 , w5592 , w5520 );
nor ( w5594 , w5593 , g12 );
nor ( w5595 , w5594 , w5340 );
not ( w5596 , w5595 );
and ( w5597 , w5596 , g11 );
not ( w5598 , w5597 );
and ( w5599 , w5598 , w5520 );
not ( w5600 , w5599 );
and ( w5601 , w5600 , w15 );
nor ( w5602 , w5587 , w5601 );
and ( w5603 , w5602 , w5520 );
and ( w5604 , w5603 , g10 );
not ( w5605 , w5604 );
and ( w5606 , w5605 , g10 );
nor ( w5607 , w5606 , w5519 );
and ( w5608 , w5744 , g4 );
and ( w5609 , w5554 , w7102 );
nor ( w5610 , w5609 , g11 );
and ( w5611 , w5610 , w5698 );
nor ( w5612 , w5611 , w4916 );
nor ( w5613 , w5608 , w5612 );
not ( w5614 , w5613 );
and ( w5615 , w5614 , w5520 );
not ( w5616 , w5147 );
and ( w5617 , w5615 , w5616 );
nor ( w5618 , w5617 , g10 );
not ( w5619 , w5618 );
and ( w5620 , w5607 , w5619 );
and ( w5621 , w5620 , w7213 );
not ( w5622 , w5621 );
and ( w5623 , w5622 , w5522 );
and ( w5624 , w5623 , w15 );
nor ( w5625 , w5624 , w4916 );
nor ( w5626 , w5583 , w5625 );
and ( w5627 , w5747 , w5520 );
and ( w5628 , w15 , w5627 );
nor ( w5629 , w5628 , w5518 );
and ( w5630 , w5629 , w5698 );
and ( w5631 , w5630 , g2 );
and ( w5632 , w5627 , g4 );
not ( w5633 , w5632 );
and ( w5634 , w5633 , w5630 );
and ( w5635 , w5634 , w7213 );
and ( w5636 , w5635 , w6380 );
nor ( w5637 , w5631 , w5636 );
nor ( w5638 , w5637 , g1 );
nor ( w5639 , w5045 , w4915 );
and ( w5640 , w5639 , w5695 );
nor ( w5641 , w5628 , w4915 );
and ( w5642 , w5640 , w5641 );
not ( w5643 , w5642 );
and ( w5644 , w5643 , w5627 );
not ( w5645 , w5644 );
and ( w5646 , w5645 , g2 );
nor ( w5647 , w5646 , w4916 );
not ( w5648 , w5627 );
and ( w5649 , w5648 , w15 );
and ( w5650 , w5647 , w5703 );
and ( w5651 , w5650 , w5627 );
nor ( w5652 , w5651 , g4 );
not ( w5653 , w5652 );
and ( w5654 , w5653 , w5520 );
nor ( w5655 , w5649 , w5519 );
and ( w5656 , w5654 , w5655 );
and ( w5657 , w5656 , g10 );
not ( w5658 , w5657 );
and ( w5659 , w5658 , g10 );
and ( w5660 , w5659 , w6380 );
not ( w5661 , w5660 );
and ( w5662 , w5627 , w5661 );
and ( w5663 , w5662 , g10 );
not ( w5664 , w5663 );
and ( w5665 , w5664 , g10 );
nor ( w5666 , w5638 , w5665 );
and ( w5667 , w5666 , w5655 );
not ( w5668 , w4916 );
and ( w5669 , w5667 , w5668 );
and ( w5670 , w5669 , g10 );
not ( w5671 , w5670 );
and ( w5672 , w5671 , g10 );
and ( w5673 , w5627 , g2 );
not ( w5674 , w5673 );
and ( w5675 , w5674 , g2 );
nor ( w5676 , w5675 , g10 );
and ( w5677 , w5676 , w5148 );
nor ( w5678 , w5677 , g10 );
nor ( w5679 , w5678 , w5340 );
not ( w5680 , w5672 );
and ( w5681 , w5680 , w5679 );
nor ( w5682 , w5681 , g12 );
nor ( w5683 , w5682 , w5340 );
not ( w5684 , w5683 );
and ( w5685 , w5684 , g11 );
and ( w5686 , w5627 , w5725 );
and ( w5687 , g11 , w5725 );
and ( w5688 , w5630 , w5765 );
and ( w5689 , w5688 , g10 );
not ( w5690 , w5689 );
and ( w5691 , w5690 , w5686 );
and ( w5692 , w5691 , w6945 );
and ( w5693 , w5686 , g10 );
nor ( w5694 , w5693 , w5687 );
not ( w5695 , w5518 );
and ( w5696 , w5694 , w5695 );
and ( w5697 , w5696 , w5752 );
not ( w5698 , w4915 );
and ( w5699 , w5697 , w5698 );
not ( w5700 , w5699 );
and ( w5701 , w5700 , g2 );
and ( w5702 , w5612 , w5725 );
not ( w5703 , w5649 );
and ( w5704 , w5702 , w5703 );
nor ( w5705 , w5704 , w5628 );
not ( w5706 , w5705 );
and ( w5707 , w5706 , g10 );
nor ( w5708 , w5707 , w4915 );
and ( w5709 , w5708 , w5765 );
and ( w5710 , w5709 , w5630 );
nor ( w5711 , w5710 , g2 );
and ( w5712 , w5711 , w7102 );
nor ( w5713 , w5701 , w5712 );
and ( w5714 , w5713 , w5765 );
not ( w5715 , w5714 );
and ( w5716 , w5715 , g1 );
and ( w5717 , w5716 , w7102 );
nor ( w5718 , w5692 , w5717 );
and ( w5719 , w5718 , w5641 );
and ( w5720 , w5719 , w5522 );
nor ( w5721 , w5720 , g4 );
nor ( w5722 , w5721 , w4915 );
and ( w5723 , w7102 , w5722 );
nor ( w5724 , w5723 , w4916 );
not ( w5725 , w5685 );
and ( w5726 , w5725 , w5724 );
and ( w5727 , w5726 , w5655 );
and ( w5728 , w5727 , g2 );
and ( w5729 , w5722 , w5641 );
and ( w5730 , w5729 , w5630 );
and ( w5731 , w5688 , w5730 );
not ( w5732 , w5728 );
and ( w5733 , w5732 , w5731 );
nor ( w5734 , w5733 , g1 );
and ( w5735 , w5731 , g2 );
not ( w5736 , w5735 );
and ( w5737 , w5736 , w5727 );
and ( w5738 , w5737 , g1 );
nor ( w5739 , w5738 , g10 );
not ( w5740 , w5734 );
and ( w5741 , w5740 , w5739 );
nor ( w5742 , w5741 , w4916 );
and ( w5743 , w5742 , w5747 );
not ( w5744 , w5519 );
and ( w5745 , w5743 , w5744 );
and ( w5746 , w5686 , w5745 );
not ( w5747 , w5626 );
and ( w5748 , w5724 , w5747 );
and ( w5749 , w5746 , w5748 );
and ( w5750 , w5749 , g2 );
nor ( w5751 , w5750 , w5518 );
not ( w5752 , w5628 );
and ( w5753 , w5751 , w5752 );
nor ( w5754 , g10 , w5741 );
not ( w5755 , w5754 );
and ( w5756 , w5755 , w5722 );
and ( w5757 , w5753 , w5756 );
not ( w5758 , w5757 );
and ( w5759 , w5758 , g1 );
nor ( w5760 , w5759 , w5687 );
nor ( w5761 , w5754 , w5518 );
and ( w5762 , w5761 , w5522 );
and ( w5763 , w5762 , w5641 );
and ( w5764 , w5763 , w5729 );
not ( w5765 , w5687 );
and ( w5766 , w5764 , w5765 );
and ( w5767 , w5760 , w5766 );
and ( w5768 , g1 , w5767 );
nor ( w5769 , w5768 , w5685 );
and ( w5770 , w5686 , w5769 );
nor ( w5771 , w5741 , w5723 );
and ( w5772 , w5770 , w5771 );
and ( w5773 , w7213 , w5772 );
nor ( w5774 , w5773 , w5518 );
and ( t_5 , w5767 , w5774 );
and ( w5775 , w6471 , g11 );
and ( w5776 , w5775 , w367 );
and ( w5777 , w5776 , w7102 );
and ( w5778 , w5777 , w15 );
nor ( w5779 , w5778 , w3 );
and ( w5780 , w2 , w5786 );
not ( w5781 , w5780 );
and ( w5782 , w5781 , w2625 );
not ( w5783 , w1735 );
and ( w5784 , w5783 , g7 );
nor ( w5785 , w5784 , w6 );
not ( w5786 , w1733 );
and ( w5787 , w5786 , w5785 );
not ( w5788 , w5787 );
and ( w5789 , w5788 , w2625 );
and ( w5790 , w5782 , w5789 );
nor ( w5791 , w5779 , w5790 );
and ( w5792 , w5791 , g10 );
and ( w5793 , w2002 , w7102 );
and ( w5794 , w5793 , w5796 );
and ( w5795 , w5794 , w5798 );
not ( w5796 , g8 );
and ( w5797 , w175 , w5796 );
not ( w5798 , g9 );
and ( w5799 , w5797 , w5798 );
and ( w5800 , w5799 , w7213 );
and ( w5801 , w5800 , w5810 );
nor ( w5802 , w5801 , w1733 );
not ( w5803 , w5802 );
and ( w5804 , w5803 , w2625 );
and ( w5805 , w5804 , w6997 );
and ( w5806 , w5805 , g11 );
nor ( w5807 , w5795 , w5806 );
not ( w5808 , w5807 );
and ( w5809 , w5808 , g13 );
not ( w5810 , w5785 );
and ( w5811 , w5809 , w5810 );
nor ( w5812 , w5811 , w1733 );
not ( w5813 , w5812 );
and ( w5814 , w5813 , w2625 );
and ( w5815 , w1796 , w7183 );
and ( w5816 , w5815 , w7213 );
and ( w5817 , w5816 , g3 );
and ( w5818 , w2333 , g11 );
nor ( w5819 , w5817 , w5818 );
nor ( w5820 , w5819 , w3 );
and ( w5821 , w5820 , w6997 );
and ( w5822 , w5821 , g11 );
nor ( w5823 , w5814 , w5822 );
nor ( w5824 , w5823 , g10 );
and ( w5825 , w5824 , g11 );
and ( w5826 , g11 , w6566 );
and ( w5827 , w5826 , g4 );
and ( w5828 , w5827 , w3 );
and ( w5829 , w5828 , w7213 );
and ( w5830 , w5829 , g3 );
and ( w5831 , w5830 , w15 );
and ( w5832 , g11 , w367 );
and ( w5833 , w5832 , w7102 );
and ( w5834 , w5833 , w3 );
and ( w5835 , w5834 , w7183 );
nor ( w5836 , w5826 , w3 );
nor ( w5837 , w5836 , w5790 );
and ( w5838 , w5837 , w7102 );
and ( w5839 , w5838 , g3 );
and ( w5840 , w5826 , w7102 );
and ( w5841 , w5840 , g2 );
and ( w5842 , w5841 , w3 );
and ( w5843 , w5842 , w6997 );
nor ( w5844 , w5839 , w5843 );
not ( w5845 , w5844 );
and ( w5846 , w5845 , w15 );
and ( w5847 , w5846 , w6997 );
nor ( w5848 , w5835 , w5847 );
nor ( w5849 , w5848 , g10 );
nor ( w5850 , w5831 , w5849 );
nor ( w5851 , w5850 , g10 );
nor ( w5852 , w5792 , w5851 );
nor ( w5853 , w92 , g11 );
nor ( w5854 , w5853 , w5822 );
nor ( w5855 , w3885 , w484 );
not ( w5856 , w5855 );
and ( w5857 , w5856 , g3 );
and ( w5858 , w5857 , w7183 );
and ( w5859 , w5854 , w5858 );
nor ( w5860 , w5859 , w3 );
nor ( w5861 , w5860 , g10 );
not ( w5862 , w5790 );
and ( w5863 , w5861 , w5862 );
and ( w5864 , w5852 , w6375 );
nor ( w5865 , w367 , g2 );
nor ( w5866 , w5865 , g2 );
nor ( w5867 , w5866 , g2 );
nor ( w5868 , w5867 , g2 );
nor ( w5869 , w5868 , w371 );
nor ( w5870 , w5869 , g1 );
and ( w5871 , w5870 , w5790 );
nor ( w5872 , w371 , w3 );
not ( w5873 , w2677 );
and ( w5874 , w5873 , w5872 );
and ( w5875 , w5874 , g3 );
nor ( w5876 , w5871 , w5875 );
not ( w5877 , w5876 );
and ( w5878 , w5877 , g3 );
not ( w5879 , w147 );
and ( w5880 , w5879 , w15 );
not ( w5881 , w5880 );
and ( w5882 , w5881 , w5790 );
and ( w5883 , w5882 , w7097 );
and ( w5884 , w15 , w5883 );
and ( w5885 , w2330 , w7183 );
and ( w5886 , w5885 , g11 );
nor ( w5887 , g13 , w5825 );
nor ( w5888 , w5887 , g3 );
and ( w5889 , w5888 , w7183 );
and ( w5890 , w5889 , w5924 );
nor ( w5891 , w5890 , g12 );
not ( w5892 , w5891 );
and ( w5893 , w5892 , w2625 );
and ( w5894 , w5893 , g11 );
nor ( w5895 , w5894 , w5825 );
and ( w5896 , w5895 , w7102 );
not ( w5897 , w5886 );
and ( w5898 , w5897 , w5896 );
nor ( w5899 , w5898 , w15 );
and ( w5900 , g13 , w5864 );
and ( w5901 , w5900 , w5924 );
not ( w5902 , w5901 );
and ( w5903 , w5902 , w15 );
nor ( w5904 , w5903 , g2 );
nor ( w5905 , w5904 , w5825 );
not ( w5906 , w5905 );
and ( w5907 , w5906 , w15 );
nor ( w5908 , w5907 , w5825 );
not ( w5909 , w5908 );
and ( w5910 , w5909 , w5790 );
and ( w5911 , w5910 , g11 );
nor ( w5912 , w5911 , w5825 );
and ( w5913 , w5912 , w7102 );
not ( w5914 , w5899 );
and ( w5915 , w5914 , w5913 );
and ( w5916 , w5915 , w6380 );
not ( w5917 , w5916 );
and ( w5918 , w5917 , w5864 );
and ( w5919 , w5918 , w2625 );
and ( w5920 , w5919 , g11 );
nor ( w5921 , w5920 , w5825 );
and ( w5922 , w5921 , w7102 );
and ( w5923 , w6049 , w5864 );
not ( w5924 , w367 );
and ( w5925 , w5923 , w5924 );
and ( w5926 , w5925 , w7183 );
and ( w5927 , w367 , w6566 );
not ( w5928 , w5927 );
and ( w5929 , w5928 , w5864 );
and ( w5930 , w5929 , w7213 );
not ( w5931 , w5930 );
and ( w5932 , w5931 , w15 );
and ( w5933 , w5932 , w6566 );
not ( w5934 , w5933 );
and ( w5935 , w5934 , w15 );
and ( w5936 , w5935 , g11 );
nor ( w5937 , w5936 , w5825 );
and ( w5938 , w5937 , w7102 );
not ( w5939 , w5926 );
and ( w5940 , w5939 , w5938 );
not ( w5941 , w5940 );
and ( w5942 , w5941 , g13 );
not ( w5943 , w5942 );
and ( w5944 , w5943 , g12 );
nor ( w5945 , w5944 , w5863 );
and ( w5946 , w5945 , w5864 );
and ( w5947 , w5946 , w5790 );
and ( w5948 , w5947 , g11 );
nor ( w5949 , w5948 , w5825 );
and ( w5950 , w5949 , w7102 );
nor ( w5951 , w5922 , w5950 );
and ( w5952 , w5951 , w2625 );
and ( w5953 , w231 , w5864 );
and ( w5954 , w5953 , w7213 );
and ( w5955 , w5954 , g3 );
and ( w5956 , w5955 , w7183 );
nor ( w5957 , w5956 , w5825 );
nor ( w5958 , w5901 , w15 );
and ( w5959 , w6471 , w367 );
nor ( w5960 , g12 , g4 );
and ( w5961 , w5960 , g13 );
not ( w5962 , w5961 );
and ( w5963 , w5962 , g11 );
not ( w5964 , w3088 );
and ( w5965 , w5964 , w5963 );
not ( w5966 , w5965 );
and ( w5967 , w5966 , g13 );
nor ( w5968 , w5967 , w3 );
and ( w5969 , w5968 , w6997 );
nor ( w5970 , w5969 , w5825 );
not ( w5971 , w5970 );
and ( w5972 , w5971 , g11 );
not ( w5973 , w5887 );
and ( w5974 , w5973 , w5972 );
and ( w5975 , w5974 , w7097 );
not ( w5976 , w5975 );
and ( w5977 , w5976 , g2 );
nor ( w5978 , w5977 , g10 );
not ( w5979 , w5959 );
and ( w5980 , w5979 , w5978 );
not ( w5981 , w5980 );
and ( w5982 , w5981 , w15 );
nor ( w5983 , w5982 , g3 );
and ( w5984 , w5983 , g11 );
nor ( w5985 , w5984 , w5825 );
and ( w5986 , w5985 , w7102 );
nor ( w5987 , w5958 , w5986 );
and ( w5988 , w5987 , w6380 );
and ( w5989 , w5900 , g2 );
and ( w5990 , w5989 , g12 );
and ( w5991 , w5990 , w6794 );
nor ( w5992 , w5991 , w5790 );
not ( w5993 , w5992 );
and ( w5994 , w5993 , g11 );
nor ( w5995 , w5865 , w5994 );
and ( w5996 , w5995 , w7183 );
and ( w5997 , g2 , w5978 );
nor ( w5998 , w1796 , w15 );
and ( w5999 , g13 , w7102 );
nor ( w6000 , w5999 , w5825 );
and ( w6001 , w6000 , w15 );
nor ( w6002 , w6001 , g3 );
and ( w6003 , w6002 , w6794 );
nor ( w6004 , w6003 , w5825 );
nor ( w6005 , w6004 , g10 );
and ( w6006 , w6005 , g11 );
not ( w6007 , w5998 );
and ( w6008 , w6007 , w6006 );
and ( w6009 , w6008 , w7097 );
and ( w6010 , w6009 , w6794 );
and ( w6011 , w6010 , w7213 );
nor ( w6012 , w6011 , w5825 );
not ( w6013 , w6012 );
and ( w6014 , g12 , w6013 );
nor ( w6015 , w5997 , w6014 );
and ( w6016 , w6015 , w15 );
nor ( w6017 , w6016 , w3 );
and ( w6018 , w6017 , g11 );
nor ( w6019 , w6018 , w5825 );
and ( w6020 , w6019 , w15 );
nor ( w6021 , w5996 , w6020 );
nor ( w6022 , w6021 , w5790 );
and ( w6023 , w6022 , w7102 );
not ( w6024 , w5988 );
and ( w6025 , w6024 , w6023 );
nor ( w6026 , w6025 , g3 );
and ( w6027 , w6026 , w6794 );
and ( w6028 , w6027 , g11 );
nor ( w6029 , w6028 , w5825 );
and ( w6030 , w6029 , w7102 );
and ( w6031 , w5957 , w6030 );
nor ( w6032 , w6031 , w3 );
and ( w6033 , w6032 , g11 );
nor ( w6034 , w6033 , w5825 );
and ( w6035 , w6034 , w7102 );
not ( w6036 , w5952 );
and ( w6037 , w6036 , w6035 );
not ( w6038 , w6037 );
and ( w6039 , g11 , w6038 );
not ( w6040 , w6039 );
and ( w6041 , g11 , w6040 );
not ( w6042 , w6041 );
and ( w6043 , w6042 , w5864 );
nor ( w6044 , w6043 , g10 );
nor ( w6045 , w401 , w6044 );
and ( w6046 , w6045 , w5789 );
and ( w6047 , w367 , w7183 );
nor ( w6048 , w6047 , g4 );
not ( w6049 , w94 );
and ( w6050 , w6049 , w6048 );
nor ( w6051 , w6050 , w5863 );
and ( w6052 , w6051 , w7183 );
and ( w6053 , w6052 , w6794 );
and ( w6054 , w367 , w7102 );
nor ( w6055 , w2002 , w6054 );
and ( w6056 , w6055 , w15 );
and ( w6057 , w6056 , w6794 );
and ( w6058 , w6057 , w7094 );
nor ( w6059 , w6058 , w6039 );
and ( w6060 , w6059 , w6997 );
not ( w6061 , w6060 );
and ( w6062 , w6061 , w5864 );
nor ( w6063 , w6062 , g10 );
and ( w6064 , w6063 , w7102 );
not ( w6065 , w6053 );
and ( w6066 , w6065 , w6064 );
nor ( w6067 , w6066 , g11 );
nor ( w6068 , w6067 , w6039 );
and ( w6069 , w6068 , w6997 );
not ( w6070 , w6046 );
and ( w6071 , w6070 , w6069 );
not ( w6072 , w6071 );
and ( w6073 , w6072 , g3 );
nor ( w6074 , w2677 , w6071 );
and ( w6075 , w6074 , w7097 );
and ( w6076 , w6075 , w5789 );
not ( w6077 , w6076 );
and ( w6078 , w6077 , w6069 );
not ( w6079 , w6073 );
and ( w6080 , w6079 , w6078 );
nor ( w6081 , w6080 , g1 );
not ( w6082 , w6081 );
and ( w6083 , w6082 , w6069 );
and ( w6084 , g7 , w5785 );
nor ( w6085 , w2002 , w6084 );
not ( w6086 , w6044 );
and ( w6087 , w6085 , w6086 );
and ( w6088 , w6087 , w5790 );
and ( w6089 , w6053 , w7094 );
nor ( w6090 , w6089 , w6039 );
and ( w6091 , w6090 , w6997 );
not ( w6092 , w6091 );
and ( w6093 , w6092 , w5864 );
nor ( w6094 , w6093 , g10 );
and ( w6095 , w6094 , w7102 );
not ( w6096 , w6088 );
and ( w6097 , w6096 , w6095 );
nor ( w6098 , w6097 , w15 );
and ( w6099 , w6098 , w6945 );
nor ( w6100 , w2002 , g4 );
and ( w6101 , w7213 , w6100 );
not ( w6102 , w6101 );
and ( w6103 , w6102 , w5789 );
not ( w6104 , w6103 );
and ( w6105 , w6104 , w6064 );
not ( w6106 , w6105 );
and ( w6107 , w6106 , w15 );
and ( w6108 , w6107 , w7094 );
nor ( w6109 , w6108 , w6039 );
and ( w6110 , w6109 , w6997 );
not ( w6111 , w6110 );
and ( w6112 , w6111 , w5864 );
nor ( w6113 , w6112 , g10 );
and ( w6114 , w6113 , w7102 );
not ( w6115 , w6099 );
and ( w6116 , w6115 , w6114 );
and ( w6117 , w6083 , w6116 );
nor ( w6118 , w6117 , g11 );
and ( w6119 , w5900 , w2625 );
and ( w6120 , w5900 , g3 );
and ( w6121 , w6120 , g2 );
and ( w6122 , w6121 , w6794 );
nor ( w6123 , w6119 , w6122 );
nor ( w6124 , w6123 , w15 );
and ( w6125 , w1904 , g3 );
nor ( w6126 , w6125 , w367 );
not ( w6127 , w231 );
and ( w6128 , w6127 , g3 );
not ( w6129 , w6128 );
and ( w6130 , w6129 , w5864 );
not ( w6131 , w6130 );
and ( w6132 , w6131 , w15 );
not ( w6133 , w6132 );
and ( w6134 , w6133 , g11 );
and ( w6135 , w6134 , w7213 );
nor ( w6136 , w6135 , w367 );
not ( w6137 , w6136 );
and ( w6138 , w6137 , w5864 );
and ( w6139 , w6138 , w15 );
and ( w6140 , w6139 , w6794 );
not ( w6141 , w6140 );
and ( w6142 , w6126 , w6141 );
not ( w6143 , w6142 );
and ( w6144 , w6143 , w5864 );
not ( w6145 , w5858 );
and ( w6146 , w6144 , w6145 );
and ( w6147 , w6146 , w15 );
and ( w6148 , w6147 , w6794 );
and ( w6149 , w6148 , g11 );
nor ( w6150 , w6149 , w5825 );
not ( w6151 , w6124 );
and ( w6152 , w6151 , w6150 );
not ( w6153 , w6152 );
and ( w6154 , w6153 , g2 );
and ( w6155 , w5864 , w5790 );
nor ( w6156 , w6155 , w5825 );
nor ( w6157 , w6156 , g13 );
and ( w6158 , w6157 , g11 );
nor ( w6159 , w234 , w6158 );
nor ( w6160 , w6159 , w15 );
not ( w6161 , w846 );
and ( w6162 , w6161 , w6150 );
not ( w6163 , w6162 );
and ( w6164 , w6163 , w15 );
and ( w6165 , w6164 , w6945 );
and ( w6166 , w2329 , w7183 );
and ( w6167 , w6166 , w5790 );
nor ( w6168 , g13 , w15 );
and ( w6169 , w2329 , w15 );
and ( w6170 , w6169 , w6794 );
and ( w6171 , w6170 , g11 );
nor ( w6172 , w6168 , w6171 );
nor ( w6173 , w6172 , w5858 );
and ( w6174 , w6173 , w6794 );
and ( w6175 , w6174 , g11 );
nor ( w6176 , w6175 , w5825 );
not ( w6177 , w6167 );
and ( w6178 , w6177 , w6176 );
and ( w6179 , w5888 , w5790 );
and ( w6180 , w2329 , w6794 );
and ( w6181 , w6180 , w7183 );
and ( w6182 , w6181 , g11 );
nor ( w6183 , w6179 , w6182 );
nor ( w6184 , w6183 , w15 );
nor ( w6185 , w6184 , w5825 );
not ( w6186 , w6185 );
and ( w6187 , w6186 , g11 );
not ( w6188 , w6187 );
and ( w6189 , w6178 , w6188 );
and ( w6190 , w6189 , g2 );
and ( w6191 , w15 , w6471 );
not ( w6192 , w6191 );
and ( w6193 , w6192 , g11 );
not ( w6194 , w527 );
and ( w6195 , w6194 , w6193 );
and ( w6196 , w6195 , w7097 );
nor ( w6197 , w6169 , w6196 );
not ( w6198 , w6197 );
and ( w6199 , w6198 , w5790 );
and ( w6200 , w5888 , g11 );
nor ( w6201 , w2329 , w6200 );
and ( w6202 , w6201 , w7183 );
not ( w6203 , w6202 );
and ( w6204 , w6203 , w6134 );
and ( w6205 , w6204 , w6794 );
nor ( w6206 , w6199 , w6205 );
and ( w6207 , w6206 , w7213 );
not ( w6208 , w6207 );
and ( w6209 , w6208 , g11 );
nor ( w6210 , w6209 , w5825 );
nor ( w6211 , w6190 , w6210 );
and ( w6212 , w6211 , g1 );
nor ( w6213 , w6212 , w5825 );
not ( w6214 , w6165 );
and ( w6215 , w6214 , w6213 );
not ( w6216 , w6215 );
and ( w6217 , w6216 , g11 );
nor ( w6218 , w6160 , w6217 );
nor ( w6219 , w6218 , w484 );
and ( w6220 , w6219 , w7213 );
and ( w6221 , w6220 , g3 );
and ( w6222 , w6471 , w5864 );
nor ( w6223 , w6222 , w15 );
nor ( w6224 , w6223 , w6191 );
and ( w6225 , w6224 , w5864 );
and ( w6226 , w6225 , w367 );
nor ( w6227 , w3891 , w6226 );
not ( w6228 , w6227 );
and ( w6229 , w6228 , w2625 );
and ( w6230 , w6222 , g2 );
and ( w6231 , w5900 , w7213 );
nor ( w6232 , w6230 , w6231 );
nor ( w6233 , w6232 , w15 );
not ( w6234 , w6233 );
and ( w6235 , w6234 , w6150 );
nor ( w6236 , w6235 , w3 );
and ( w6237 , w6236 , g11 );
nor ( w6238 , w6229 , w6237 );
nor ( w6239 , w6238 , w5858 );
and ( w6240 , w6239 , w7097 );
and ( w6241 , w6240 , w6945 );
not ( w6242 , w6241 );
and ( w6243 , w6242 , w6213 );
not ( w6244 , w6243 );
and ( w6245 , w6244 , g10 );
and ( w6246 , w6039 , w6997 );
nor ( w6247 , w6245 , w6246 );
not ( w6248 , w6247 );
and ( w6249 , w6248 , g11 );
nor ( w6250 , w6249 , g4 );
not ( w6251 , w6221 );
and ( w6252 , w6251 , w6250 );
nor ( w6253 , w6252 , g1 );
not ( w6254 , w6253 );
and ( w6255 , w6254 , w6213 );
not ( w6256 , w6255 );
and ( w6257 , w6256 , g10 );
nor ( w6258 , w6257 , w6246 );
not ( w6259 , w6258 );
and ( w6260 , w6259 , g11 );
nor ( w6261 , w6260 , g4 );
not ( w6262 , w6154 );
and ( w6263 , w6262 , w6261 );
not ( w6264 , w6263 );
and ( w6265 , w6264 , g3 );
not ( w6266 , w6265 );
and ( w6267 , w6266 , w6250 );
nor ( w6268 , w6267 , g1 );
not ( w6269 , w6268 );
and ( w6270 , w6269 , w6213 );
not ( w6271 , w6270 );
and ( w6272 , w6271 , g10 );
nor ( w6273 , w6272 , w6246 );
not ( w6274 , w6273 );
and ( w6275 , w6274 , g11 );
and ( w6276 , w6275 , w5864 );
nor ( w6277 , w6276 , g4 );
not ( w6278 , w6118 );
and ( w6279 , w6278 , w6277 );
not ( w6280 , w6279 );
and ( w6281 , w15 , w6280 );
and ( w6282 , w6281 , w6794 );
not ( w6283 , w6282 );
and ( w6284 , w6283 , g10 );
nor ( w6285 , w6284 , w6117 );
not ( w6286 , w6285 );
and ( w6287 , w6286 , w6277 );
not ( w6288 , w5884 );
and ( w6289 , w6288 , w6287 );
nor ( w6290 , w5789 , w150 );
not ( w6291 , w6290 );
and ( w6292 , w6291 , g2 );
not ( w6293 , w6292 );
and ( w6294 , w6293 , g10 );
nor ( w6295 , w6294 , w6117 );
and ( w6296 , w6295 , w7094 );
not ( w6297 , w6296 );
and ( w6298 , w6297 , w6277 );
and ( w6299 , w6289 , w6298 );
nor ( w6300 , w6299 , g3 );
not ( w6301 , w6300 );
and ( w6302 , w6301 , g10 );
nor ( w6303 , w6302 , w6117 );
and ( w6304 , w6303 , w7094 );
not ( w6305 , w6304 );
and ( w6306 , w6305 , w6277 );
not ( w6307 , w5878 );
and ( w6308 , w6307 , w6306 );
and ( w6309 , w6308 , g10 );
nor ( w6310 , w6309 , w6117 );
and ( w6311 , w6310 , w7094 );
not ( w6312 , w6311 );
and ( w6313 , w6312 , w6277 );
and ( w6314 , w5864 , w6942 );
and ( w6315 , w6314 , g13 );
nor ( w6316 , g4 , w6313 );
and ( w6317 , w6896 , g10 );
nor ( w6318 , w6317 , w6313 );
and ( w6319 , w6318 , g13 );
nor ( w6320 , w3437 , w6316 );
not ( w6321 , w6320 );
and ( w6322 , w6321 , g11 );
nor ( w6323 , w6316 , w6322 );
nor ( w6324 , w6323 , w6313 );
and ( w6325 , w6324 , w6945 );
nor ( w6326 , w6325 , w6316 );
nor ( w6327 , g13 , w6313 );
nor ( w6328 , w6327 , w6316 );
nor ( w6329 , w6328 , w15 );
nor ( w6330 , w6316 , g13 );
nor ( w6331 , w6330 , w6313 );
and ( w6332 , w15 , w6331 );
nor ( w6333 , w6332 , w6316 );
not ( w6334 , w6333 );
and ( w6335 , w6334 , g3 );
nor ( w6336 , w6335 , w6316 );
not ( w6337 , w6329 );
and ( w6338 , w6337 , w6336 );
nor ( w6339 , w6338 , g10 );
and ( w6340 , w6339 , g3 );
nor ( w6341 , w6340 , w6316 );
not ( w6342 , w6341 );
and ( w6343 , w6342 , g11 );
nor ( w6344 , w6316 , w6343 );
not ( w6345 , w6330 );
and ( w6346 , w6345 , g10 );
nor ( w6347 , w6346 , w6316 );
nor ( w6348 , w6347 , w6313 );
nor ( w6349 , w6348 , w15 );
nor ( w6350 , w5997 , w6316 );
and ( w6351 , w6350 , w6566 );
and ( w6352 , w6896 , g2 );
nor ( w6353 , w6331 , g2 );
nor ( w6354 , w6353 , w6313 );
not ( w6355 , w6352 );
and ( w6356 , w6355 , w6354 );
and ( w6357 , w6356 , g10 );
nor ( w6358 , w6357 , w6316 );
nor ( w6359 , w6358 , w3 );
and ( w6360 , w6359 , g11 );
nor ( w6361 , w6360 , w6316 );
and ( w6362 , w6361 , w6566 );
and ( w6363 , w6351 , w6362 );
and ( w6364 , w6363 , w15 );
nor ( w6365 , w6364 , w6313 );
and ( w6366 , w6365 , w6794 );
and ( w6367 , w7097 , w6366 );
not ( w6368 , w6349 );
and ( w6369 , w6368 , w6367 );
nor ( w6370 , w6369 , w6316 );
and ( w6371 , w6370 , g2 );
not ( w6372 , w6331 );
and ( w6373 , w6372 , g10 );
nor ( w6374 , w6373 , w6313 );
not ( w6375 , w5863 );
and ( w6376 , w6374 , w6375 );
and ( w6377 , w6376 , g3 );
nor ( w6378 , w6200 , w6316 );
nor ( w6379 , w6378 , w6313 );
not ( w6380 , g12 );
and ( w6381 , g13 , w6380 );
and ( w6382 , w527 , w6794 );
and ( w6383 , w6382 , w6997 );
nor ( w6384 , w6381 , w6383 );
nor ( w6385 , w6384 , w15 );
and ( w6386 , w6385 , w6945 );
and ( w6387 , w15 , w5978 );
and ( w6388 , w6387 , w6794 );
and ( w6389 , w6388 , w7097 );
nor ( w6390 , w6386 , w6389 );
nor ( w6391 , w527 , w6389 );
not ( w6392 , w6391 );
and ( w6393 , w6392 , g1 );
and ( w6394 , w6393 , w6794 );
and ( w6395 , w6394 , w6997 );
nor ( w6396 , w6395 , w5825 );
and ( w6397 , w6390 , w6396 );
nor ( w6398 , w6397 , w3 );
and ( w6399 , w6398 , w6997 );
and ( w6400 , w6379 , w6399 );
nor ( w6401 , w6400 , w6316 );
and ( w6402 , w6401 , w6566 );
not ( w6403 , w6377 );
and ( w6404 , w6403 , w6402 );
nor ( w6405 , w6404 , w15 );
and ( w6406 , w6331 , g3 );
nor ( w6407 , w6406 , w6367 );
and ( w6408 , w6407 , w6896 );
not ( w6409 , w6408 );
and ( w6410 , w6409 , g10 );
nor ( w6411 , w6410 , w6316 );
not ( w6412 , w6411 );
and ( w6413 , w6412 , w15 );
nor ( w6414 , w6413 , w6316 );
nor ( w6415 , w6414 , w3 );
and ( w6416 , w6415 , g11 );
nor ( w6417 , w6416 , w6316 );
and ( w6418 , w6417 , w6566 );
not ( w6419 , w6405 );
and ( w6420 , w6419 , w6418 );
and ( w6421 , w3097 , w5864 );
nor ( w6422 , w6421 , w6316 );
nor ( w6423 , w6422 , w6313 );
nor ( w6424 , w6423 , w5825 );
nor ( w6425 , w6424 , g10 );
nor ( w6426 , w6425 , w6316 );
not ( w6427 , w6426 );
and ( w6428 , w6427 , g3 );
nor ( w6429 , w6316 , w15 );
not ( w6430 , w6429 );
and ( w6431 , w6430 , w6366 );
nor ( w6432 , w6431 , w6316 );
nor ( w6433 , w6432 , g3 );
nor ( w6434 , w6433 , w6316 );
not ( w6435 , w6428 );
and ( w6436 , w6435 , w6434 );
nor ( w6437 , w6436 , w3 );
and ( w6438 , w6437 , g11 );
not ( w6439 , w6438 );
and ( w6440 , w6420 , w6439 );
and ( w6441 , w6440 , w7213 );
nor ( w6442 , w6441 , w6313 );
and ( w6443 , w6442 , w6794 );
and ( w6444 , w6443 , g11 );
not ( w6445 , w6371 );
and ( w6446 , w6445 , w6444 );
nor ( w6447 , w6446 , w6316 );
and ( w6448 , w6447 , w6566 );
and ( w6449 , w6344 , w6448 );
and ( w6450 , w6449 , g2 );
not ( w6451 , w6450 );
and ( w6452 , w6451 , w6444 );
nor ( w6453 , w6452 , w6316 );
not ( w6454 , w6453 );
and ( w6455 , w6454 , g1 );
nor ( w6456 , w6455 , w6316 );
and ( w6457 , w6456 , w6566 );
and ( w6458 , w6326 , w6457 );
nor ( w6459 , w6458 , w3 );
and ( w6460 , w6459 , w7213 );
nor ( w6461 , w6460 , w6316 );
nor ( w6462 , w6461 , g10 );
nor ( w6463 , w6462 , w6316 );
not ( w6464 , w6463 );
and ( w6465 , w6464 , w15 );
nor ( w6466 , w6465 , w6316 );
not ( w6467 , w6466 );
and ( w6468 , w6467 , g3 );
nor ( w6469 , w6468 , w6316 );
and ( w6470 , w6469 , w6566 );
not ( w6471 , g13 );
and ( w6472 , w6471 , w6470 );
and ( w6473 , w6472 , g1 );
not ( w6474 , w6473 );
and ( w6475 , w6474 , g11 );
and ( w6476 , w6475 , g13 );
and ( w6477 , w6379 , w2625 );
and ( w6478 , w6222 , w6942 );
nor ( w6479 , w6478 , w6316 );
nor ( w6480 , w6479 , g1 );
and ( w6481 , w6480 , w7097 );
nor ( w6482 , w6481 , w6316 );
and ( w6483 , w6482 , w6457 );
nor ( w6484 , w6483 , w3 );
and ( w6485 , w6484 , g2 );
and ( w6486 , w6896 , g13 );
not ( w6487 , w6486 );
and ( w6488 , w6487 , w5864 );
nor ( w6489 , w6488 , g1 );
nor ( w6490 , w230 , w6313 );
and ( w6491 , w6490 , g11 );
not ( w6492 , w6489 );
and ( w6493 , w6492 , w6491 );
nor ( w6494 , w6493 , w6316 );
not ( w6495 , w6494 );
and ( w6496 , w6495 , g3 );
and ( w6497 , w6496 , w2625 );
nor ( w6498 , w6497 , w6316 );
nor ( w6499 , w5900 , w6316 );
not ( w6500 , w6499 );
and ( w6501 , w6500 , g3 );
nor ( w6502 , w6330 , g3 );
and ( w6503 , w6502 , w6945 );
not ( w6504 , w6503 );
and ( w6505 , w6504 , w6457 );
nor ( w6506 , w6505 , w3 );
nor ( w6507 , w6506 , w6316 );
not ( w6508 , w6507 );
and ( w6509 , w6508 , g10 );
nor ( w6510 , w6509 , w6316 );
and ( w6511 , w6331 , w6945 );
nor ( w6512 , w6511 , w6316 );
and ( w6513 , w6512 , w6457 );
nor ( w6514 , w6513 , w3 );
nor ( w6515 , w6514 , w6316 );
not ( w6516 , w6515 );
and ( w6517 , w6516 , g2 );
nor ( w6518 , w6517 , w6316 );
not ( w6519 , w6518 );
and ( w6520 , w6519 , g3 );
nor ( w6521 , w6520 , w6316 );
not ( w6522 , w6521 );
and ( w6523 , w6522 , w15 );
and ( w6524 , w6523 , g11 );
nor ( w6525 , w6524 , w6316 );
and ( w6526 , w6331 , w2625 );
nor ( w6527 , w6526 , w6316 );
not ( w6528 , w5978 );
and ( w6529 , w6527 , w6528 );
nor ( w6530 , w6529 , w6313 );
and ( w6531 , w6530 , g2 );
nor ( w6532 , w6531 , w6316 );
nor ( w6533 , w6532 , g3 );
nor ( w6534 , w6533 , w5825 );
not ( w6535 , w2 );
and ( w6536 , w6535 , g2 );
and ( w6537 , w6536 , g4 );
nor ( w6538 , w6537 , w5825 );
nor ( w6539 , w6538 , w5785 );
nor ( w6540 , w6539 , w1733 );
not ( w6541 , w6540 );
and ( w6542 , w6541 , w2625 );
nor ( w6543 , w6542 , w6389 );
not ( w6544 , w6543 );
and ( w6545 , w15 , w6544 );
nor ( w6546 , w6545 , w5825 );
nor ( w6547 , w6546 , g10 );
not ( w6548 , w6534 );
and ( w6549 , w6548 , w6547 );
nor ( w6550 , w6549 , w6316 );
not ( w6551 , w6550 );
and ( w6552 , w15 , w6551 );
nor ( w6553 , w6552 , w6316 );
and ( w6554 , w6553 , w6470 );
not ( w6555 , w6554 );
and ( w6556 , w6555 , g11 );
nor ( w6557 , w6556 , w6316 );
and ( w6558 , w6525 , w6557 );
nor ( w6559 , w6558 , g10 );
nor ( w6560 , w6559 , w6316 );
and ( w6561 , w6510 , w6560 );
not ( w6562 , w6561 );
and ( w6563 , w6562 , w15 );
and ( w6564 , w6563 , g11 );
nor ( w6565 , w6564 , w6316 );
not ( w6566 , w5825 );
and ( w6567 , w6565 , w6566 );
not ( w6568 , w6501 );
and ( w6569 , w6568 , w6567 );
nor ( w6570 , w6313 , w5863 );
not ( w6571 , w6569 );
and ( w6572 , w6571 , w6570 );
and ( w6573 , w6572 , w6945 );
nor ( w6574 , w6573 , w6316 );
and ( w6575 , w6574 , w6457 );
nor ( w6576 , w6575 , w3 );
nor ( w6577 , w6576 , w6316 );
nor ( w6578 , w6577 , g2 );
nor ( w6579 , w6578 , w6316 );
not ( w6580 , w6579 );
and ( w6581 , w6580 , g10 );
nor ( w6582 , w6581 , w6316 );
and ( w6583 , w6582 , w6560 );
not ( w6584 , w6583 );
and ( w6585 , w15 , w6584 );
nor ( w6586 , w6585 , w6316 );
and ( w6587 , w6586 , w6470 );
not ( w6588 , w6587 );
and ( w6589 , w6588 , g11 );
nor ( w6590 , w6589 , w6316 );
and ( w6591 , w6498 , w6590 );
nor ( w6592 , w6591 , g2 );
nor ( w6593 , w6592 , w6316 );
not ( w6594 , w6593 );
and ( w6595 , w6594 , g10 );
nor ( w6596 , w6595 , w6316 );
and ( w6597 , w6596 , w6560 );
not ( w6598 , w6597 );
and ( w6599 , w15 , w6598 );
nor ( w6600 , w6599 , w6316 );
and ( w6601 , w6600 , w6470 );
not ( w6602 , w6485 );
and ( w6603 , w6602 , w6601 );
not ( w6604 , w6603 );
and ( w6605 , w6604 , g10 );
not ( w6606 , w6605 );
and ( w6607 , w6606 , w6560 );
not ( w6608 , w6607 );
and ( w6609 , w15 , w6608 );
nor ( w6610 , w6609 , w6316 );
and ( w6611 , w6610 , w6470 );
not ( w6612 , w6611 );
and ( w6613 , w6612 , g11 );
nor ( w6614 , w6477 , w6613 );
and ( w6615 , w6614 , w6896 );
not ( w6616 , w6615 );
and ( w6617 , w6616 , g2 );
nor ( w6618 , w6617 , w6316 );
and ( w6619 , w6618 , w6601 );
not ( w6620 , w6619 );
and ( w6621 , w6620 , g10 );
nor ( w6622 , w6621 , w6316 );
and ( w6623 , w6622 , w6560 );
not ( w6624 , w6623 );
and ( w6625 , w15 , w6624 );
nor ( w6626 , w6625 , w6316 );
and ( w6627 , w6626 , w6470 );
not ( w6628 , w6476 );
and ( w6629 , w6628 , w6627 );
not ( w6630 , w6629 );
and ( w6631 , w6630 , w6570 );
and ( w6632 , w6631 , w7097 );
and ( w6633 , w6632 , g10 );
nor ( w6634 , w6633 , w6316 );
nor ( w6635 , w6634 , g2 );
nor ( w6636 , w6635 , w6316 );
not ( w6637 , w6636 );
and ( w6638 , w6637 , w5790 );
nor ( w6639 , w6638 , w6316 );
and ( w6640 , w6222 , w6997 );
nor ( w6641 , w6640 , w6316 );
nor ( w6642 , w6641 , w6313 );
and ( w6643 , w6642 , g2 );
nor ( w6644 , w6643 , w6316 );
not ( w6645 , w6373 );
and ( w6646 , w6645 , w5864 );
and ( w6647 , w6646 , w6942 );
and ( w6648 , w6647 , w7213 );
nor ( w6649 , w6648 , w6316 );
and ( w6650 , w6644 , w6649 );
not ( w6651 , w6650 );
and ( w6652 , w6651 , g3 );
and ( w6653 , w6331 , g2 );
and ( w6654 , w6653 , g10 );
nor ( w6655 , w6654 , w6316 );
nor ( w6656 , w6655 , g3 );
nor ( w6657 , w6656 , w6316 );
nor ( w6658 , w6657 , w15 );
nor ( w6659 , w6652 , w6658 );
nor ( w6660 , w6659 , g1 );
nor ( w6661 , w6660 , w6316 );
and ( w6662 , w6661 , w6457 );
nor ( w6663 , w6662 , w3 );
nor ( w6664 , w6663 , w6316 );
nor ( w6665 , w6664 , w15 );
nor ( w6666 , w6665 , w6316 );
and ( w6667 , w6666 , w6627 );
not ( w6668 , w6667 );
and ( w6669 , w6668 , g11 );
nor ( w6670 , w6669 , w6316 );
and ( w6671 , w6639 , w6670 );
nor ( w6672 , w6671 , w15 );
nor ( w6673 , w6672 , w6316 );
and ( w6674 , w6673 , w6627 );
not ( w6675 , w6319 );
and ( w6676 , w6675 , w6674 );
not ( w6677 , w6676 );
and ( w6678 , w6677 , g3 );
nor ( w6679 , w6678 , w6316 );
not ( w6680 , w6679 );
and ( w6681 , w6680 , g2 );
not ( w6682 , w6681 );
and ( w6683 , w6682 , w6674 );
not ( w6684 , w6683 );
and ( w6685 , w6684 , w5789 );
nor ( w6686 , w6685 , w6316 );
and ( w6687 , w6686 , w6670 );
nor ( w6688 , w6687 , w15 );
nor ( w6689 , w6688 , w6316 );
and ( w6690 , w6689 , w6627 );
not ( w6691 , w6690 );
and ( w6692 , w6691 , g11 );
nor ( w6693 , w6692 , w6316 );
not ( w6694 , w6315 );
and ( w6695 , w6694 , w6693 );
not ( w6696 , w6695 );
and ( w6697 , w6696 , w2625 );
nor ( w6698 , w6697 , w6316 );
nor ( w6699 , w6698 , g2 );
nor ( w6700 , w6699 , w6316 );
not ( w6701 , w6700 );
and ( w6702 , w6701 , g3 );
nor ( w6703 , w6702 , w6316 );
not ( w6704 , w6703 );
and ( w6705 , w6704 , g10 );
nor ( w6706 , w6705 , w6316 );
not ( w6707 , w6084 );
and ( w6708 , w2625 , w6707 );
and ( w6709 , w6708 , w5790 );
and ( w6710 , w6457 , w6627 );
not ( w6711 , w6709 );
and ( w6712 , w6711 , w6710 );
nor ( w6713 , w6712 , w6313 );
and ( w6714 , w6713 , g2 );
nor ( w6715 , w578 , w6014 );
and ( w6716 , w6715 , w6457 );
nor ( w6717 , w6716 , w3 );
nor ( w6718 , w6717 , w6316 );
nor ( w6719 , w6718 , w6313 );
and ( w6720 , w6719 , w6997 );
nor ( w6721 , w6720 , w6316 );
nor ( w6722 , w6721 , w15 );
nor ( w6723 , w6722 , w6316 );
and ( w6724 , w6723 , w6627 );
not ( w6725 , w6724 );
and ( w6726 , w6725 , g11 );
nor ( w6727 , w6726 , w6316 );
nor ( w6728 , w6727 , g2 );
nor ( w6729 , w6728 , w6316 );
nor ( w6730 , w6729 , g10 );
nor ( w6731 , w6730 , w6316 );
and ( w6732 , w6731 , w6693 );
not ( w6733 , w6714 );
and ( w6734 , w6733 , w6732 );
not ( w6735 , w6734 );
and ( w6736 , w6735 , g13 );
not ( w6737 , w6736 );
and ( w6738 , w6737 , w6693 );
nor ( w6739 , w6738 , g3 );
nor ( w6740 , w6739 , w6316 );
nor ( w6741 , w6740 , g10 );
nor ( w6742 , w6741 , w6316 );
and ( w6743 , w6742 , w6693 );
nor ( w6744 , w6743 , w15 );
not ( w6745 , w6744 );
and ( w6746 , w6745 , w6627 );
not ( w6747 , w6746 );
and ( w6748 , w6747 , g11 );
nor ( w6749 , w6748 , w6316 );
and ( w6750 , w6703 , w6749 );
nor ( w6751 , w6750 , g10 );
nor ( w6752 , w6751 , w6316 );
and ( w6753 , w6752 , w6693 );
nor ( w6754 , w6753 , w15 );
nor ( w6755 , w6754 , w6316 );
and ( w6756 , w6755 , w6627 );
not ( w6757 , w6756 );
and ( w6758 , w6757 , g11 );
nor ( w6759 , w6758 , w6316 );
and ( w6760 , w6706 , w6759 );
nor ( w6761 , w6760 , w15 );
nor ( w6762 , w6761 , w6316 );
and ( w6763 , w6762 , w6627 );
not ( w6764 , w6763 );
and ( w6765 , w6764 , g11 );
nor ( w6766 , w6765 , w6316 );
and ( w6767 , g11 , w6766 );
nor ( w6768 , w6767 , w6313 );
and ( w6769 , w6768 , w5789 );
and ( w6770 , w6965 , g1 );
and ( w6771 , w6770 , w6942 );
not ( w6772 , w6771 );
and ( w6773 , w6772 , w6766 );
nor ( w6774 , w6773 , w3 );
nor ( w6775 , w6774 , w6316 );
not ( w6776 , w6769 );
and ( w6777 , w6776 , w6775 );
nor ( w6778 , w15 , w6777 );
not ( w6779 , w6778 );
and ( w6780 , w6779 , w6766 );
not ( w6781 , w6780 );
and ( w6782 , w6781 , g10 );
and ( w6783 , w6766 , w7183 );
and ( w6784 , w6783 , w3 );
not ( w6785 , w6784 );
and ( w6786 , w6785 , w5864 );
and ( w6787 , w6786 , w6570 );
and ( w6788 , w6787 , w6965 );
and ( w6789 , w6788 , w6945 );
not ( w6790 , w6783 );
and ( w6791 , w6790 , w5864 );
and ( w6792 , w6791 , w5790 );
and ( w6793 , w6570 , w7183 );
not ( w6794 , w3 );
and ( w6795 , w6793 , w6794 );
nor ( w6796 , w6792 , w6795 );
and ( w6797 , w6796 , w6766 );
nor ( w6798 , w6797 , g10 );
nor ( w6799 , w6789 , w6798 );
and ( w6800 , w6799 , w6896 );
and ( w6801 , w6800 , w6997 );
nor ( w6802 , w6801 , g10 );
nor ( w6803 , w6802 , w6316 );
not ( w6804 , w6803 );
and ( w6805 , w6804 , g3 );
nor ( w6806 , w6805 , w6316 );
not ( w6807 , w6782 );
and ( w6808 , w6807 , w6806 );
nor ( w6809 , w6808 , w6313 );
and ( w6810 , w6809 , g3 );
not ( w6811 , w6788 );
and ( w6812 , w6811 , g10 );
nor ( w6813 , w6783 , w6313 );
and ( w6814 , w6813 , w6965 );
and ( w6815 , w6814 , w5790 );
not ( w6816 , w6815 );
and ( w6817 , w6816 , w6766 );
and ( w6818 , w6817 , w6997 );
nor ( w6819 , w6818 , w6767 );
and ( w6820 , w6819 , w6945 );
nor ( w6821 , w6820 , w6316 );
nor ( w6822 , w6821 , g3 );
nor ( w6823 , w6822 , w6316 );
nor ( w6824 , w6812 , w6823 );
and ( w6825 , w6824 , w6945 );
and ( w6826 , w6814 , g10 );
not ( w6827 , w6826 );
and ( w6828 , w6827 , w6766 );
and ( w6829 , w6828 , w3 );
and ( w6830 , w6768 , g10 );
and ( w6831 , w6623 , w15 );
nor ( w6832 , w6831 , w6313 );
and ( w6833 , w6832 , w6965 );
and ( w6834 , w6833 , w6997 );
and ( w6835 , w6834 , g1 );
nor ( w6836 , w6830 , w6835 );
not ( w6837 , w6836 );
and ( w6838 , w6837 , g1 );
not ( w6839 , w6829 );
and ( w6840 , w6839 , w6838 );
nor ( w6841 , w6825 , w6840 );
nor ( w6842 , w6841 , g3 );
nor ( w6843 , w6842 , w6316 );
not ( w6844 , w6810 );
and ( w6845 , w6844 , w6843 );
and ( w6846 , w6845 , w7213 );
nor ( w6847 , w6846 , w6313 );
and ( w6848 , w6965 , w6847 );
and ( w6849 , w6848 , g3 );
nor ( w6850 , w6846 , g2 );
and ( w6851 , w6766 , w6855 );
and ( w6852 , w6848 , w7183 );
not ( w6853 , w6852 );
and ( w6854 , w6853 , w6766 );
not ( w6855 , w6850 );
and ( w6856 , w6854 , w6855 );
not ( w6857 , w6856 );
and ( w6858 , w6857 , g3 );
and ( w6859 , w6851 , w7183 );
nor ( w6860 , w6859 , w6313 );
and ( w6861 , w6860 , w6965 );
and ( w6862 , w6861 , w6847 );
and ( w6863 , w6862 , w7097 );
nor ( w6864 , w6863 , w6850 );
not ( w6865 , w6864 );
and ( w6866 , w6865 , g1 );
and ( w6867 , w6866 , g10 );
nor ( w6868 , w6858 , w6867 );
not ( w6869 , w6868 );
and ( w6870 , w6869 , g10 );
not ( w6871 , w6870 );
and ( w6872 , w6851 , w6871 );
not ( w6873 , w6872 );
and ( w6874 , w6873 , g10 );
nor ( w6875 , w6773 , w6846 );
nor ( w6876 , w6875 , w6850 );
not ( w6877 , w6876 );
and ( w6878 , w6877 , g3 );
nor ( w6879 , w6862 , g10 );
nor ( w6880 , w6879 , g10 );
nor ( w6881 , w6850 , w6316 );
not ( w6882 , w6880 );
and ( w6883 , w6882 , w6881 );
nor ( w6884 , w6883 , w3 );
nor ( w6885 , w6884 , w6316 );
and ( w6886 , w6885 , w6881 );
not ( w6887 , w6878 );
and ( w6888 , w6887 , w6886 );
and ( w6889 , w6888 , w7183 );
not ( w6890 , w6889 );
and ( w6891 , w6890 , w6848 );
and ( w6892 , w6891 , w6997 );
nor ( w6893 , w6892 , w6316 );
nor ( w6894 , w6893 , w3 );
nor ( w6895 , w6874 , w6894 );
not ( w6896 , w6316 );
and ( w6897 , w6895 , w6896 );
nor ( w6898 , w6897 , w3 );
nor ( w6899 , w6898 , w6316 );
and ( w6900 , w6899 , w6881 );
not ( w6901 , w6849 );
and ( w6902 , w6901 , w6900 );
nor ( w6903 , w6902 , g1 );
nor ( w6904 , w6903 , w6870 );
not ( w6905 , w6904 );
and ( w6906 , w6905 , g10 );
nor ( w6907 , w6906 , w6894 );
nor ( w6908 , w6907 , w3 );
nor ( w6909 , w5789 , w6908 );
nor ( w6910 , w6909 , w6846 );
nor ( w6911 , w6909 , w6313 );
and ( w6912 , w6910 , w6911 );
and ( w6913 , w6848 , w6912 );
and ( w6914 , w6913 , w7183 );
not ( w6915 , w6908 );
and ( w6916 , w6851 , w6915 );
not ( w6917 , w6914 );
and ( w6918 , w6917 , w6916 );
not ( w6919 , w6918 );
and ( w6920 , w6919 , g3 );
and ( w6921 , w15 , w6916 );
nor ( w6922 , w6921 , w6909 );
and ( w6923 , w6922 , w6965 );
and ( w6924 , w6923 , w6945 );
not ( w6925 , w6924 );
and ( w6926 , w6925 , w6916 );
nor ( w6927 , w6926 , w6313 );
not ( w6928 , w6846 );
and ( w6929 , w6927 , w6928 );
and ( w6930 , w6929 , w7097 );
nor ( w6931 , w6930 , g10 );
nor ( w6932 , w6931 , g10 );
nor ( w6933 , w6920 , w6932 );
and ( w6934 , w6933 , w6997 );
nor ( w6935 , w6934 , g10 );
nor ( w6936 , w6935 , w6850 );
nor ( w6937 , w6908 , w6850 );
and ( w6938 , w6936 , w6937 );
nor ( w6939 , w6767 , w6909 );
not ( w6940 , w6934 );
and ( w6941 , w6939 , w6940 );
not ( w6942 , w6313 );
and ( w6943 , w6941 , w6942 );
and ( w6944 , w6943 , w7183 );
not ( w6945 , g1 );
and ( w6946 , w6766 , w6945 );
nor ( w6947 , w6946 , w6767 );
nor ( w6948 , w6934 , w6313 );
and ( w6949 , w6948 , w6847 );
and ( w6950 , w6949 , w6912 );
and ( w6951 , w6947 , w6950 );
not ( w6952 , w6951 );
and ( w6953 , w6952 , w6881 );
nor ( w6954 , w6935 , w6316 );
and ( w6955 , w6954 , w6937 );
and ( w6956 , w6953 , w6955 );
not ( w6957 , w6956 );
and ( w6958 , w6957 , w15 );
nor ( w6959 , w6944 , w6958 );
nor ( w6960 , w6959 , w6846 );
and ( w6961 , w6960 , w7097 );
nor ( w6962 , g3 , w6961 );
nor ( w6963 , w6962 , w6313 );
and ( w6964 , w6963 , w6950 );
not ( w6965 , w6767 );
and ( w6966 , w6964 , w6965 );
and ( w6967 , w15 , w6966 );
nor ( w6968 , w6967 , w6908 );
and ( w6969 , w6968 , w6937 );
and ( w6970 , w6938 , w6969 );
not ( w6971 , w6961 );
and ( w6972 , w6970 , w6971 );
nand ( t_6 , w6972 , w6766 );
not ( w6973 , w92 );
and ( w6974 , w15 , w6973 );
and ( w6975 , w2292 , w15 );
not ( w6976 , w6975 );
and ( w6977 , w6976 , g3 );
nor ( w6978 , w374 , g3 );
and ( w6979 , w6978 , w7094 );
nor ( w6980 , w6977 , w6979 );
and ( w6981 , w6980 , g4 );
nor ( w6982 , w457 , g3 );
and ( w6983 , w6982 , w7094 );
not ( w6984 , w6983 );
and ( w6985 , g2 , w6984 );
nor ( w6986 , w6985 , g3 );
nor ( w6987 , w94 , w6986 );
and ( w6988 , w6987 , w7183 );
and ( w6989 , w6988 , w7102 );
nor ( w6990 , w6989 , g11 );
not ( w6991 , w6981 );
and ( w6992 , w6991 , w6990 );
and ( w6993 , w1746 , w7183 );
nor ( w6994 , w6993 , w494 );
and ( w6995 , w6994 , g3 );
nor ( w6996 , w6995 , w6983 );
not ( w6997 , g10 );
and ( w6998 , w6996 , w6997 );
nor ( w6999 , w6998 , g11 );
not ( w7000 , w6999 );
and ( w7001 , w7000 , w228 );
not ( w7002 , w7001 );
and ( w7003 , w6992 , w7002 );
not ( w7004 , w7003 );
and ( w7005 , w7004 , w228 );
and ( w7006 , w6974 , w7060 );
not ( w7007 , w7006 );
and ( w7008 , w7007 , g10 );
nor ( w7009 , w7005 , w15 );
nor ( w7010 , w7009 , g10 );
not ( w7011 , w7010 );
and ( w7012 , w7011 , g3 );
and ( w7013 , w7060 , g10 );
nor ( w7014 , w7013 , g2 );
and ( w7015 , w7014 , g4 );
nor ( w7016 , w7015 , w7005 );
and ( w7017 , w7016 , w7183 );
and ( w7018 , g11 , w228 );
nor ( w7019 , w7018 , g2 );
nor ( w7020 , w7019 , g10 );
nor ( w7021 , w7020 , w7005 );
and ( w7022 , w7021 , g4 );
not ( w7023 , w7018 );
and ( w7024 , w7023 , g2 );
and ( w7025 , w7013 , w7213 );
and ( w7026 , w7025 , w7102 );
and ( w7027 , w15 , w7026 );
and ( w7028 , w7027 , w7097 );
and ( w7029 , w7028 , w7094 );
not ( w7030 , w7029 );
and ( w7031 , w7030 , w228 );
not ( w7032 , w7024 );
and ( w7033 , w7032 , w7031 );
nor ( w7034 , w7033 , g4 );
and ( w7035 , w15 , w7034 );
and ( w7036 , w7035 , w7097 );
and ( w7037 , w7036 , w7094 );
not ( w7038 , w7037 );
and ( w7039 , w7038 , w228 );
not ( w7040 , w7022 );
and ( w7041 , w7040 , w7039 );
not ( w7042 , w7041 );
and ( w7043 , w15 , w7042 );
and ( w7044 , w7043 , w7097 );
and ( w7045 , w7044 , w7094 );
not ( w7046 , w7045 );
and ( w7047 , w7046 , w228 );
not ( w7048 , w7017 );
and ( w7049 , w7048 , w7047 );
nor ( w7050 , w7049 , g3 );
and ( w7051 , w7050 , w7094 );
not ( w7052 , w7051 );
and ( w7053 , w7052 , w228 );
not ( w7054 , w7012 );
and ( w7055 , w7054 , w7053 );
nor ( w7056 , w7055 , g11 );
not ( w7057 , w7056 );
and ( w7058 , w7057 , w228 );
nor ( w7059 , g2 , w7058 );
not ( w7060 , w7005 );
and ( w7061 , w7060 , g2 );
and ( w7062 , w7061 , w15 );
and ( w7063 , w7062 , g3 );
not ( w7064 , w7063 );
and ( w7065 , w7064 , w7053 );
not ( w7066 , w7059 );
and ( w7067 , w7066 , w7065 );
and ( w7068 , w7067 , g4 );
nor ( w7069 , w7009 , g4 );
not ( w7070 , w7069 );
and ( w7071 , w7070 , g3 );
not ( w7072 , w7071 );
and ( w7073 , w7072 , w7053 );
nor ( w7074 , w7073 , g11 );
not ( w7075 , w7074 );
and ( w7076 , w7075 , w228 );
nor ( w7077 , w7068 , w7076 );
nor ( w7078 , w7077 , g10 );
not ( w7079 , w7078 );
and ( w7080 , w7079 , g3 );
not ( w7081 , w7080 );
and ( w7082 , w7081 , w7053 );
nor ( w7083 , w7008 , w7082 );
and ( w7084 , w7083 , g3 );
not ( w7085 , w7084 );
and ( w7086 , w7085 , w7053 );
and ( w7087 , w7213 , w7086 );
nor ( w7088 , w7087 , w15 );
not ( w7089 , w7088 );
and ( w7090 , w7089 , w7086 );
nor ( w7091 , w7090 , w7005 );
not ( w7092 , w7082 );
and ( w7093 , w7091 , w7092 );
not ( w7094 , g11 );
and ( w7095 , w7093 , w7094 );
and ( w7096 , w7095 , w7213 );
not ( w7097 , g3 );
and ( w7098 , w7096 , w7097 );
nor ( w7099 , w7098 , g4 );
not ( w7100 , w7099 );
and ( w7101 , w7100 , w7093 );
not ( w7102 , g4 );
and ( w7103 , w7101 , w7102 );
not ( w7104 , g7 );
and ( w7105 , w7104 , w7093 );
not ( w7106 , w11 );
and ( w7107 , w7106 , w7093 );
and ( w7108 , w7105 , w7107 );
nor ( w7109 , w7103 , w7108 );
nor ( w7110 , w1733 , w7108 );
not ( w7111 , w7110 );
and ( w7112 , w7111 , w7107 );
and ( w7113 , w7109 , w7205 );
and ( w7114 , w7113 , g2 );
not ( w7115 , w7114 );
and ( w7116 , w7115 , w7095 );
and ( w7117 , w7116 , w7183 );
and ( w7118 , w7095 , g10 );
not ( w7119 , w7118 );
and ( w7120 , w7119 , w7113 );
nor ( w7121 , w7120 , g2 );
not ( w7122 , w7121 );
and ( w7123 , w7122 , g4 );
and ( w7124 , w7095 , g2 );
nor ( w7125 , w7124 , w7101 );
nor ( w7126 , w7125 , g3 );
not ( w7127 , w7123 );
and ( w7128 , w7127 , w7126 );
not ( w7129 , w7128 );
and ( w7130 , w7113 , w7129 );
not ( w7131 , w7130 );
and ( w7132 , w7131 , w15 );
nor ( w7133 , w7132 , w7112 );
and ( w7134 , w7133 , w7113 );
not ( w7135 , w7134 );
and ( w7136 , w7135 , g10 );
nor ( w7137 , w7136 , w7112 );
and ( w7138 , w7113 , w7183 );
not ( w7139 , w7095 );
and ( w7140 , w15 , w7139 );
not ( w7141 , w7140 );
and ( w7142 , w7141 , w7093 );
not ( w7143 , w7138 );
and ( w7144 , w7143 , w7142 );
and ( w7145 , w7144 , g2 );
and ( w7146 , w7095 , w7183 );
and ( w7147 , w7133 , g4 );
not ( w7148 , w7147 );
and ( w7149 , w7148 , w7126 );
nor ( w7150 , w7146 , w7149 );
nor ( w7151 , w7150 , g2 );
not ( w7152 , w7151 );
and ( w7153 , w7152 , g4 );
not ( w7154 , w7153 );
and ( w7155 , w7154 , w7126 );
nor ( w7156 , w7145 , w7155 );
nor ( w7157 , w7156 , g10 );
not ( w7158 , w7157 );
and ( w7159 , w7158 , g4 );
not ( w7160 , w7159 );
and ( w7161 , w7160 , w7126 );
and ( w7162 , w7137 , w7170 );
and ( w7163 , w7162 , g4 );
not ( w7164 , w7163 );
and ( w7165 , w7164 , w7126 );
nor ( w7166 , w7117 , w7165 );
not ( w7167 , w7166 );
and ( w7168 , w7167 , g10 );
nor ( w7169 , w7168 , w7112 );
not ( w7170 , w7161 );
and ( w7171 , w7169 , w7170 );
and ( w7172 , w7171 , g4 );
not ( w7173 , w7172 );
and ( w7174 , w7173 , w7126 );
and ( w7175 , w7113 , w7207 );
and ( w7176 , w7175 , g2 );
nor ( w7177 , g3 , w7174 );
and ( w7178 , g11 , w7109 );
nor ( w7179 , w7177 , w7178 );
and ( w7180 , w7095 , w7179 );
not ( w7181 , w7176 );
and ( w7182 , w7181 , w7180 );
not ( w7183 , w15 );
and ( w7184 , w7182 , w7183 );
and ( w7185 , w7175 , g10 );
not ( w7186 , w7185 );
and ( w7187 , w7186 , w7180 );
not ( w7188 , w7187 );
and ( w7189 , w7188 , g2 );
not ( w7190 , w7180 );
and ( w7191 , w15 , w7190 );
not ( w7192 , w7191 );
and ( w7193 , w7192 , w7093 );
and ( w7194 , w7228 , w7093 );
and ( w7195 , w7193 , w7194 );
not ( w7196 , w7189 );
and ( w7197 , w7196 , w7195 );
and ( w7198 , w7197 , w7180 );
and ( w7199 , w15 , w7198 );
nor ( w7200 , w7199 , w7112 );
and ( w7201 , w7200 , w7113 );
and ( w7202 , w7201 , w7207 );
nor ( w7203 , w7202 , g4 );
nor ( w7204 , w7184 , w7203 );
not ( w7205 , w7112 );
and ( w7206 , w7204 , w7205 );
not ( w7207 , w7174 );
and ( w7208 , w7206 , w7207 );
nor ( w7209 , w7208 , g4 );
nor ( w7210 , w7209 , w7112 );
nor ( w7211 , w7209 , w7174 );
and ( w7212 , w7210 , w7211 );
not ( w7213 , g2 );
and ( w7214 , w7212 , w7213 );
and ( w7215 , w7214 , w15 );
nor ( w7216 , w7215 , w7177 );
and ( w7217 , w7216 , w7093 );
not ( w7218 , w7217 );
and ( w7219 , w7218 , g10 );
not ( w7220 , w7219 );
and ( w7221 , w7220 , w7093 );
not ( w7222 , w7214 );
and ( w7223 , w7222 , w7093 );
nor ( w7224 , w7223 , w15 );
and ( w7225 , w7212 , g2 );
nor ( w7226 , g4 , w7209 );
nor ( w7227 , w7225 , w7226 );
not ( w7228 , w7177 );
and ( w7229 , w7227 , w7228 );
not ( w7230 , w7229 );
and ( w7231 , w7230 , w15 );
nor ( w7232 , w7224 , w7231 );
nor ( w7233 , w7232 , g10 );
not ( w7234 , w7233 );
and ( w7235 , w7234 , w7180 );
and ( w7236 , w7221 , w7235 );
nor ( w7237 , w7226 , w7177 );
and ( w7238 , w7237 , w7180 );
and ( t_7 , w7236 , w7238 );

endmodule
