module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 ; 
output g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 ; 
wire t_0 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( g157 , n158 ); 
buf ( g158 , n159 ); 
buf ( g159 , n160 ); 
buf ( g160 , n161 ); 
buf ( g161 , n162 ); 
buf ( g162 , n163 ); 
buf ( g163 , n164 ); 
buf ( g164 , n165 ); 
buf ( g165 , n166 ); 
buf ( g166 , n167 ); 
buf ( g167 , n168 ); 
buf ( g168 , n169 ); 
buf ( g169 , n170 ); 
buf ( g170 , n171 ); 
buf ( g171 , n172 ); 
buf ( g172 , n173 ); 
buf ( g173 , n174 ); 
buf ( g174 , n175 ); 
buf ( g175 , n176 ); 
buf ( g176 , n177 ); 
buf ( g177 , n178 ); 
buf ( g178 , n179 ); 
buf ( g179 , n180 ); 
buf ( g180 , n181 ); 
buf ( g181 , n182 ); 
buf ( g182 , n183 ); 
buf ( g183 , n184 ); 
buf ( g184 , n185 ); 
buf ( g185 , n186 ); 
buf ( g186 , n187 ); 
buf ( g187 , n188 ); 
buf ( g188 , n189 ); 
buf ( g189 , n190 ); 
buf ( g190 , n191 ); 
buf ( g191 , n192 ); 
buf ( g192 , n193 ); 
buf ( g193 , n194 ); 
buf ( g194 , n195 ); 
buf ( g195 , n196 ); 
buf ( g196 , n197 ); 
buf ( g197 , n198 ); 
buf ( g198 , n199 ); 
buf ( g199 , n200 ); 
buf ( g200 , n201 ); 
buf ( g201 , n202 ); 
buf ( g202 , n203 ); 
buf ( g203 , n204 ); 
buf ( g204 , n205 ); 
buf ( g205 , n206 ); 
buf ( g206 , n207 ); 
buf ( g207 , n208 ); 
buf ( g208 , n209 ); 
buf ( g209 , n210 ); 
buf ( g210 , n211 ); 
buf ( g211 , n212 ); 
buf ( g212 , n213 ); 
buf ( g213 , n214 ); 
buf ( g214 , n215 ); 
buf ( g215 , n216 ); 
buf ( g216 , n217 ); 
buf ( g217 , n218 ); 
buf ( g218 , n219 ); 
buf ( g219 , n220 ); 
buf ( g220 , n221 ); 
buf ( n158 , n115 ); 
buf ( n159 , n115 ); 
buf ( n160 , n115 ); 
buf ( n161 , n124 ); 
buf ( n162 , n124 ); 
buf ( n163 , n137 ); 
buf ( n164 , n137 ); 
buf ( n165 , n137 ); 
buf ( n166 , n1056 ); 
buf ( n167 , n1053 ); 
buf ( n168 , n1060 ); 
buf ( n169 , n1055 ); 
buf ( n170 , n1059 ); 
buf ( n171 , n1057 ); 
buf ( n172 , n1058 ); 
buf ( n173 , n1054 ); 
buf ( n174 , n1049 ); 
buf ( n175 , n1048 ); 
buf ( n176 , n115 ); 
buf ( n177 , n1052 ); 
buf ( n178 , n1042 ); 
buf ( n179 , n1044 ); 
buf ( n180 , n1046 ); 
buf ( n181 , n1040 ); 
buf ( n182 , n1041 ); 
buf ( n183 , n593 ); 
buf ( n184 , n477 ); 
buf ( n185 , n1037 ); 
buf ( n186 , n747 ); 
buf ( n187 , n770 ); 
buf ( n188 , n1031 ); 
buf ( n189 , n373 ); 
buf ( n190 , n1035 ); 
buf ( n191 , n1036 ); 
buf ( n192 , n1039 ); 
buf ( n193 , n244 ); 
buf ( n194 , n378 ); 
buf ( n195 , n1034 ); 
buf ( n196 , n400 ); 
buf ( n197 , n348 ); 
buf ( n198 , n448 ); 
buf ( n199 , n494 ); 
buf ( n200 , n1029 ); 
buf ( n201 , n1029 ); 
buf ( n202 , n1033 ); 
buf ( n203 , n1033 ); 
buf ( n204 , n1023 ); 
buf ( n205 , n1026 ); 
buf ( n206 , n1026 ); 
buf ( n207 , n1020 ); 
buf ( n208 , n675 ); 
buf ( n209 , n651 ); 
buf ( n210 , n628 ); 
buf ( n211 , n976 ); 
buf ( n212 , n977 ); 
buf ( n213 , n1017 ); 
buf ( n214 , n1001 ); 
buf ( n215 , n1000 ); 
buf ( n216 , n1000 ); 
buf ( n217 , n1002 ); 
buf ( n218 , n588 ); 
buf ( n219 , 1'b0 ); 
buf ( n220 , n837 ); 
buf ( n221 , n838 ); 
not ( n229 , n49 ); 
not ( n230 , n117 ); 
nand ( n231 , n230 , n120 ); 
not ( n232 , n231 ); 
not ( n233 , n232 ); 
or ( n234 , n229 , n233 ); 
nand ( n235 , n120 , n60 , n117 ); 
nand ( n236 , n234 , n235 ); 
not ( n237 , n236 ); 
not ( n238 , n120 ); 
and ( n239 , n117 , n39 ); 
not ( n240 , n117 ); 
and ( n241 , n240 , n71 ); 
or ( n242 , n239 , n241 ); 
nand ( n243 , n238 , n242 ); 
nand ( n244 , n237 , n243 ); 
not ( n245 , n244 ); 
not ( n246 , n146 ); 
not ( n247 , n246 ); 
not ( n248 , n110 ); 
nor ( n249 , n248 , n145 ); 
not ( n250 , n249 ); 
or ( n251 , n247 , n250 ); 
nand ( n252 , n146 , n90 , n145 ); 
nand ( n253 , n251 , n252 ); 
not ( n254 , n145 ); 
nand ( n255 , n254 , n146 , n100 ); 
not ( n256 , n146 ); 
nand ( n257 , n256 , n80 , n145 ); 
nand ( n258 , n255 , n257 ); 
nor ( n259 , n253 , n258 ); 
not ( n260 , n259 ); 
not ( n261 , n146 ); 
nand ( n262 , n261 , n79 , n145 ); 
not ( n263 , n145 ); 
nand ( n264 , n263 , n146 , n99 ); 
nand ( n265 , n262 , n264 ); 
not ( n266 , n146 ); 
not ( n267 , n109 ); 
nor ( n268 , n267 , n145 ); 
nand ( n269 , n266 , n268 ); 
nand ( n270 , n146 , n89 , n145 ); 
nand ( n271 , n269 , n270 ); 
nor ( n272 , n265 , n271 ); 
not ( n273 , n127 ); 
and ( n274 , n260 , n272 , n273 , n30 ); 
buf ( n275 , n274 ); 
and ( n276 , n275 , n139 ); 
not ( n277 , n275 ); 
and ( n278 , n277 , n128 ); 
nor ( n279 , n276 , n278 ); 
not ( n280 , n279 ); 
or ( n281 , n245 , n280 ); 
or ( n282 , n244 , n279 ); 
nand ( n283 , n281 , n282 ); 
and ( n284 , n275 , n138 ); 
not ( n285 , n275 ); 
and ( n286 , n285 , n126 ); 
nor ( n287 , n284 , n286 ); 
nand ( n288 , n61 , n117 ); 
and ( n289 , n120 , n288 ); 
not ( n290 , n120 ); 
not ( n291 , n117 ); 
nand ( n292 , n291 , n72 ); 
and ( n293 , n290 , n292 ); 
or ( n294 , n289 , n293 ); 
not ( n295 , n120 ); 
nand ( n296 , n295 , n40 , n117 ); 
not ( n297 , n231 ); 
nand ( n298 , n50 , n297 ); 
nand ( n299 , n294 , n296 , n298 ); 
not ( n300 , n299 ); 
not ( n301 , n300 ); 
not ( n302 , n301 ); 
not ( n303 , n302 ); 
not ( n304 , n303 ); 
nand ( n305 , n283 , n287 , n304 ); 
not ( n306 , n243 ); 
nor ( n307 , n236 , n306 ); 
nand ( n308 , n307 , n279 ); 
not ( n309 , n42 ); 
not ( n310 , n231 ); 
not ( n311 , n310 ); 
or ( n312 , n309 , n311 ); 
not ( n313 , n120 ); 
nand ( n314 , n313 , n31 , n117 ); 
nand ( n315 , n312 , n314 ); 
nand ( n316 , n120 , n52 , n117 ); 
not ( n317 , n120 ); 
not ( n318 , n117 ); 
nand ( n319 , n317 , n63 , n318 ); 
nand ( n320 , n316 , n319 ); 
nor ( n321 , n315 , n320 ); 
not ( n322 , n136 ); 
not ( n323 , n303 ); 
not ( n324 , n287 ); 
or ( n325 , n323 , n324 ); 
or ( n326 , n303 , n287 ); 
nand ( n327 , n325 , n326 ); 
nand ( n328 , t_0 , n327 , n283 ); 
nand ( n329 , n305 , n308 , n328 ); 
nor ( n330 , n259 , n127 ); 
and ( n331 , n330 , n272 , n30 ); 
not ( n332 , n331 ); 
not ( n333 , n132 ); 
nand ( n334 , n332 , n333 , n8 ); 
not ( n335 , n334 ); 
not ( n336 , n335 ); 
not ( n337 , n275 ); 
nand ( n338 , n120 , n318 ); 
not ( n339 , n338 ); 
not ( n340 , n339 ); 
nand ( n341 , n120 , n56 , n117 ); 
not ( n342 , n120 ); 
nand ( n343 , n342 , n35 , n117 ); 
not ( n344 , n120 ); 
nand ( n345 , n344 , n67 , n318 ); 
nand ( n346 , n340 , n341 , n343 , n345 ); 
not ( n347 , n346 ); 
not ( n348 , n347 ); 
nand ( n349 , n337 , n8 , n348 ); 
not ( n350 , n349 ); 
not ( n351 , n350 ); 
or ( n352 , n336 , n351 ); 
nand ( n353 , n334 , n349 ); 
nand ( n354 , n352 , n353 ); 
not ( n355 , n275 ); 
or ( n356 , n140 , n355 ); 
not ( n357 , n129 ); 
not ( n358 , n275 ); 
nand ( n359 , n357 , n358 ); 
nand ( n360 , n356 , n359 ); 
nand ( n361 , n59 , n117 ); 
and ( n362 , n120 , n361 ); 
not ( n363 , n120 ); 
nand ( n364 , n38 , n117 ); 
and ( n365 , n363 , n364 ); 
nor ( n366 , n362 , n365 ); 
not ( n367 , n48 ); 
not ( n368 , n297 ); 
or ( n369 , n367 , n368 ); 
not ( n370 , n120 ); 
nand ( n371 , n370 , n70 , n318 ); 
nand ( n372 , n369 , n371 ); 
nor ( n373 , n366 , n372 ); 
and ( n374 , n360 , n373 ); 
not ( n375 , n360 ); 
not ( n376 , n366 ); 
nand ( n377 , n48 , n339 ); 
nand ( n378 , n376 , n377 , n371 ); 
and ( n379 , n375 , n378 ); 
nor ( n380 , n374 , n379 ); 
not ( n381 , n131 ); 
nor ( n382 , n381 , n331 ); 
not ( n383 , n142 ); 
not ( n384 , n331 ); 
or ( n385 , n383 , n384 ); 
nand ( n386 , n385 , n8 ); 
nor ( n387 , n382 , n386 ); 
not ( n388 , n46 ); 
not ( n389 , n338 ); 
not ( n390 , n389 ); 
or ( n391 , n388 , n390 ); 
not ( n392 , n120 ); 
nand ( n393 , n392 , n36 , n117 ); 
nand ( n394 , n391 , n393 ); 
not ( n395 , n394 ); 
nand ( n396 , n120 , n57 , n117 ); 
not ( n397 , n120 ); 
nand ( n398 , n397 , n68 , n318 ); 
and ( n399 , n396 , n398 ); 
nand ( n400 , n395 , n399 ); 
nand ( n401 , n8 , n400 ); 
not ( n402 , n401 ); 
and ( n403 , n387 , n402 ); 
not ( n404 , n387 ); 
and ( n405 , n404 , n401 ); 
nor ( n406 , n403 , n405 ); 
not ( n407 , n406 ); 
nand ( n408 , n354 , n380 , n407 ); 
not ( n409 , n141 ); 
not ( n410 , n331 ); 
or ( n411 , n409 , n410 ); 
nand ( n412 , n411 , n8 ); 
not ( n413 , n130 ); 
nor ( n414 , n413 , n331 ); 
nor ( n415 , n412 , n414 ); 
and ( n416 , n120 , n58 , n117 ); 
not ( n417 , n69 ); 
nor ( n418 , n417 , n120 , n117 ); 
nor ( n419 , n416 , n418 ); 
nand ( n420 , n37 , n117 ); 
nor ( n421 , n120 , n420 ); 
not ( n422 , n421 ); 
nand ( n423 , n47 , n339 ); 
nand ( n424 , n419 , n422 , n423 ); 
nand ( n425 , n8 , n424 ); 
and ( n426 , n415 , n425 ); 
not ( n427 , n415 ); 
not ( n428 , n425 ); 
and ( n429 , n427 , n428 ); 
nor ( n430 , n426 , n429 ); 
not ( n431 , n331 ); 
not ( n432 , n133 ); 
nand ( n433 , n431 , n432 , n8 ); 
not ( n434 , n433 ); 
not ( n435 , n275 ); 
and ( n436 , n45 , n232 ); 
nand ( n437 , n34 , n117 ); 
nor ( n438 , n120 , n437 ); 
nor ( n439 , n436 , n438 ); 
nand ( n440 , n55 , n117 ); 
not ( n441 , n440 ); 
and ( n442 , n120 , n441 ); 
not ( n443 , n120 ); 
not ( n444 , n66 ); 
nor ( n445 , n444 , n117 ); 
and ( n446 , n443 , n445 ); 
nor ( n447 , n442 , n446 ); 
nand ( n448 , n439 , n447 ); 
nand ( n449 , n435 , n8 , n448 ); 
xor ( n450 , n434 , n449 ); 
nand ( n451 , n430 , n450 ); 
nor ( n452 , n408 , n451 ); 
and ( n453 , n329 , n452 ); 
nand ( n454 , n407 , n430 ); 
nand ( n455 , n373 , n360 ); 
nand ( n456 , n354 , n450 ); 
nor ( n457 , n454 , n455 , n456 ); 
nor ( n458 , n453 , n457 ); 
and ( n459 , n450 , n335 , n349 ); 
and ( n460 , n434 , n449 ); 
nor ( n461 , n459 , n460 ); 
not ( n462 , n461 ); 
nand ( n463 , n415 , n450 ); 
not ( n464 , n406 ); 
nand ( n465 , n464 , n354 , n425 ); 
nor ( n466 , n463 , n465 ); 
buf ( n467 , n387 ); 
nand ( n468 , n354 , n467 ); 
nand ( n469 , n401 , n450 ); 
nor ( n470 , n468 , n469 ); 
nor ( n471 , n462 , n466 , n470 ); 
nand ( n472 , n458 , n471 ); 
not ( n473 , n134 ); 
not ( n474 , n330 ); 
nor ( n475 , n265 , n271 ); 
not ( n476 , n475 ); 
not ( n477 , n476 ); 
nand ( n478 , n474 , n477 , n30 ); 
not ( n479 , n478 ); 
not ( n480 , n275 ); 
and ( n481 , n473 , n479 , n480 ); 
not ( n482 , n481 ); 
nand ( n483 , n54 , n117 ); 
not ( n484 , n483 ); 
and ( n485 , n120 , n484 ); 
not ( n486 , n120 ); 
not ( n487 , n65 ); 
nor ( n488 , n487 , n117 ); 
and ( n489 , n486 , n488 ); 
nor ( n490 , n485 , n489 ); 
not ( n491 , n120 ); 
nand ( n492 , n491 , n33 , n117 ); 
nand ( n493 , n44 , n339 ); 
nand ( n494 , n490 , n492 , n493 ); 
and ( n495 , n494 , n479 , n480 ); 
not ( n496 , n495 ); 
or ( n497 , n482 , n496 ); 
or ( n498 , n481 , n495 ); 
nand ( n499 , n497 , n498 ); 
not ( n500 , n135 ); 
and ( n501 , n500 , n479 , n355 ); 
not ( n502 , n275 ); 
not ( n503 , n95 ); 
not ( n504 , n146 ); 
nor ( n505 , n504 , n145 ); 
not ( n506 , n505 ); 
or ( n507 , n503 , n506 ); 
nand ( n508 , n145 , n146 ); 
not ( n509 , n508 ); 
nand ( n510 , n85 , n509 ); 
nand ( n511 , n507 , n510 ); 
not ( n512 , n75 ); 
not ( n513 , n145 ); 
nor ( n514 , n513 , n146 ); 
not ( n515 , n514 ); 
or ( n516 , n512 , n515 ); 
nor ( n517 , n145 , n146 ); 
nand ( n518 , n105 , n517 ); 
nand ( n519 , n516 , n518 ); 
nor ( n520 , n511 , n519 ); 
not ( n521 , n520 ); 
nand ( n522 , n502 , n521 , n479 ); 
xor ( n523 , n501 , n522 ); 
not ( n524 , n275 ); 
not ( n525 , n138 ); 
nand ( n526 , n524 , n525 , n479 ); 
not ( n527 , n526 ); 
not ( n528 , n527 ); 
not ( n529 , n275 ); 
not ( n530 , n92 ); 
not ( n531 , n530 ); 
nand ( n532 , n145 , n146 ); 
not ( n533 , n532 ); 
and ( n534 , n531 , n533 ); 
nor ( n535 , n145 , n146 ); 
and ( n536 , n112 , n535 ); 
nor ( n537 , n534 , n536 ); 
not ( n538 , n146 ); 
nor ( n539 , n538 , n145 ); 
nand ( n540 , n102 , n539 ); 
not ( n541 , n145 ); 
nor ( n542 , n541 , n146 ); 
nand ( n543 , n82 , n542 ); 
nand ( n544 , n537 , n540 , n543 ); 
not ( n545 , n544 ); 
not ( n546 , n545 ); 
nand ( n547 , n529 , n546 , n479 ); 
not ( n548 , n547 ); 
not ( n549 , n548 ); 
or ( n550 , n528 , n549 ); 
nand ( n551 , n526 , n547 ); 
nand ( n552 , n550 , n551 ); 
not ( n553 , n275 ); 
nand ( n554 , n553 , n322 , n479 ); 
not ( n555 , n554 ); 
not ( n556 , n555 ); 
and ( n557 , n103 , n539 ); 
not ( n558 , n93 ); 
nor ( n559 , n558 , n532 ); 
nor ( n560 , n557 , n559 ); 
and ( n561 , n83 , n542 ); 
and ( n562 , n113 , n517 ); 
nor ( n563 , n561 , n562 ); 
nand ( n564 , n560 , n563 ); 
and ( n565 , n564 , n479 , n355 ); 
not ( n566 , n565 ); 
or ( n567 , n556 , n566 ); 
or ( n568 , n555 , n565 ); 
nand ( n569 , n567 , n568 ); 
and ( n570 , n499 , n523 , n552 , n569 ); 
not ( n571 , n565 ); 
nand ( n572 , n552 , n571 , n555 ); 
and ( n573 , n501 , n522 ); 
nand ( n574 , n573 , n552 , n569 ); 
and ( n575 , n572 , n574 ); 
nand ( n576 , n527 , n547 ); 
nand ( n577 , n481 , n552 , n523 ); 
not ( n578 , n577 ); 
not ( n579 , n569 ); 
nor ( n580 , n579 , n495 ); 
nand ( n581 , n578 , n580 ); 
nand ( n582 , n575 , n576 , n581 ); 
nor ( n583 , n570 , n582 ); 
and ( n584 , n472 , n583 ); 
not ( n585 , n472 ); 
not ( n586 , n582 ); 
and ( n587 , n585 , n586 ); 
nor ( n588 , n584 , n587 ); 
nand ( n589 , n32 , n76 , n64 , n106 ); 
and ( n590 , n147 , n589 ); 
nand ( n591 , n53 , n86 , n43 , n96 ); 
and ( n592 , n119 , n591 ); 
nor ( n593 , n590 , n592 ); 
or ( n594 , n500 , n136 ); 
or ( n595 , n322 , n135 ); 
nand ( n596 , n594 , n595 ); 
not ( n597 , n596 ); 
and ( n598 , n133 , n473 ); 
and ( n599 , n134 , n432 ); 
nor ( n600 , n598 , n599 ); 
not ( n601 , n600 ); 
or ( n602 , n597 , n601 ); 
or ( n603 , n600 , n596 ); 
nand ( n604 , n602 , n603 ); 
not ( n605 , n604 ); 
and ( n606 , n129 , n413 ); 
not ( n607 , n129 ); 
and ( n608 , n607 , n130 ); 
nor ( n609 , n606 , n608 ); 
not ( n610 , n156 ); 
not ( n611 , n128 ); 
not ( n612 , n611 ); 
or ( n613 , n610 , n612 ); 
not ( n614 , n156 ); 
nand ( n615 , n614 , n128 ); 
nand ( n616 , n613 , n615 ); 
and ( n617 , n131 , n132 ); 
not ( n618 , n131 ); 
and ( n619 , n618 , n333 ); 
nor ( n620 , n617 , n619 ); 
xor ( n621 , n616 , n620 ); 
and ( n622 , n609 , n621 ); 
nor ( n623 , n609 , n621 ); 
nor ( n624 , n622 , n623 ); 
not ( n625 , n624 ); 
and ( n626 , n605 , n625 ); 
and ( n627 , n604 , n624 ); 
nor ( n628 , n626 , n627 ); 
not ( n629 , n628 ); 
nand ( n630 , n593 , n629 ); 
xor ( n631 , n143 , n144 ); 
not ( n632 , n631 ); 
not ( n633 , n139 ); 
and ( n634 , n140 , n633 ); 
not ( n635 , n140 ); 
and ( n636 , n635 , n139 ); 
nor ( n637 , n634 , n636 ); 
xor ( n638 , n138 , n157 ); 
and ( n639 , n141 , n142 ); 
not ( n640 , n141 ); 
not ( n641 , n142 ); 
and ( n642 , n640 , n641 ); 
nor ( n643 , n639 , n642 ); 
xor ( n644 , n638 , n643 ); 
and ( n645 , n637 , n644 ); 
nor ( n646 , n637 , n644 ); 
nor ( n647 , n645 , n646 ); 
not ( n648 , n647 ); 
and ( n649 , n632 , n648 ); 
and ( n650 , n631 , n647 ); 
nor ( n651 , n649 , n650 ); 
xor ( n652 , n154 , n155 ); 
not ( n653 , n126 ); 
and ( n654 , n125 , n653 ); 
not ( n655 , n125 ); 
and ( n656 , n655 , n126 ); 
nor ( n657 , n654 , n656 ); 
xnor ( n658 , n652 , n657 ); 
and ( n659 , n148 , n149 ); 
not ( n660 , n148 ); 
not ( n661 , n149 ); 
and ( n662 , n660 , n661 ); 
nor ( n663 , n659 , n662 ); 
and ( n664 , n152 , n153 ); 
not ( n665 , n152 ); 
not ( n666 , n153 ); 
and ( n667 , n665 , n666 ); 
nor ( n668 , n664 , n667 ); 
xor ( n669 , n663 , n668 ); 
xnor ( n670 , n150 , n151 ); 
xor ( n671 , n669 , n670 ); 
and ( n672 , n658 , n671 ); 
or ( n673 , n658 , n671 ); 
nand ( n674 , n673 , n10 ); 
nor ( n675 , n672 , n674 ); 
nor ( n676 , n651 , n675 ); 
not ( n677 , n97 ); 
not ( n678 , n505 ); 
or ( n679 , n677 , n678 ); 
not ( n680 , n532 ); 
nand ( n681 , n87 , n680 ); 
nand ( n682 , n679 , n681 ); 
not ( n683 , n77 ); 
not ( n684 , n514 ); 
or ( n685 , n683 , n684 ); 
nand ( n686 , n107 , n535 ); 
nand ( n687 , n685 , n686 ); 
nor ( n688 , n682 , n687 ); 
and ( n689 , 1'b1 , n688 ); 
nor ( n690 , n689 , 1'b0 ); 
not ( n691 , n690 ); 
and ( n692 , n146 , n88 ); 
not ( n693 , n146 ); 
and ( n694 , n693 , n78 ); 
or ( n695 , n692 , n694 ); 
nand ( n696 , n695 , n145 ); 
not ( n697 , n145 ); 
and ( n698 , n146 , n98 ); 
not ( n699 , n146 ); 
and ( n700 , n699 , n108 ); 
or ( n701 , n698 , n700 ); 
nand ( n702 , n697 , n701 ); 
nand ( n703 , n696 , n702 ); 
and ( n704 , n703 , n476 ); 
not ( n705 , n703 ); 
and ( n706 , n705 , n477 ); 
nor ( n707 , n704 , n706 ); 
not ( n708 , n707 ); 
and ( n709 , n691 , n708 ); 
and ( n710 , n690 , n707 ); 
nor ( n711 , n709 , n710 ); 
not ( n712 , n711 ); 
not ( n713 , n712 ); 
not ( n714 , n94 ); 
not ( n715 , n714 ); 
not ( n716 , n508 ); 
and ( n717 , n715 , n716 ); 
and ( n718 , n114 , n535 ); 
nor ( n719 , n717 , n718 ); 
nand ( n720 , n104 , n505 ); 
nand ( n721 , n84 , n514 ); 
nand ( n722 , n719 , n720 , n721 ); 
not ( n723 , n722 ); 
not ( n724 , n520 ); 
or ( n725 , n723 , n724 ); 
not ( n726 , n722 ); 
nand ( n727 , n521 , n726 ); 
nand ( n728 , n725 , n727 ); 
not ( n729 , n728 ); 
and ( n730 , n81 , n542 ); 
not ( n731 , n91 ); 
nor ( n732 , n731 , n532 ); 
nor ( n733 , n730 , n732 ); 
and ( n734 , n101 , n539 ); 
and ( n735 , n111 , n517 ); 
nor ( n736 , n734 , n735 ); 
nand ( n737 , n733 , n736 ); 
not ( n738 , n252 ); 
not ( n739 , n110 ); 
nor ( n740 , n739 , n146 , n145 ); 
nor ( n741 , n738 , n740 ); 
buf ( n742 , n257 ); 
buf ( n743 , n255 ); 
nand ( n744 , n741 , n742 , n743 ); 
and ( n745 , n737 , n744 ); 
not ( n746 , n737 ); 
not ( n747 , n744 ); 
and ( n748 , n746 , n747 ); 
nor ( n749 , n745 , n748 ); 
not ( n750 , n749 ); 
or ( n751 , n729 , n750 ); 
or ( n752 , n728 , n749 ); 
nand ( n753 , n751 , n752 ); 
and ( n754 , n564 , n545 ); 
not ( n755 , n564 ); 
and ( n756 , n755 , n546 ); 
nor ( n757 , n754 , n756 ); 
and ( n758 , n753 , n757 ); 
not ( n759 , n753 ); 
not ( n760 , n757 ); 
and ( n761 , n759 , n760 ); 
nor ( n762 , n758 , n761 ); 
not ( n763 , n762 ); 
not ( n764 , n763 ); 
or ( n765 , n713 , n764 ); 
and ( n766 , n711 , n762 ); 
nor ( n767 , n766 , n29 ); 
nand ( n768 , n765 , n767 ); 
not ( n769 , n399 ); 
nor ( n770 , n394 , n769 ); 
xor ( n771 , n770 , n347 ); 
not ( n772 , n771 ); 
not ( n773 , n772 ); 
not ( n774 , n494 ); 
and ( n775 , n448 , n774 ); 
not ( n776 , n448 ); 
and ( n777 , n776 , n494 ); 
nor ( n778 , n775 , n777 ); 
not ( n779 , n778 ); 
not ( n780 , n779 ); 
or ( n781 , n773 , n780 ); 
nand ( n782 , n771 , n778 ); 
nand ( n783 , n781 , n782 ); 
not ( n784 , n783 ); 
not ( n785 , n784 ); 
and ( n786 , n47 , n389 ); 
nor ( n787 , n786 , n421 ); 
nand ( n788 , n787 , n419 ); 
and ( n789 , n788 , n378 ); 
not ( n790 , n788 ); 
and ( n791 , n790 , n373 ); 
nor ( n792 , n789 , n791 ); 
not ( n793 , n792 ); 
not ( n794 , n320 ); 
nand ( n795 , n42 , n389 ); 
nand ( n796 , n794 , n314 , n795 ); 
not ( n797 , n796 ); 
nand ( n798 , n62 , n117 ); 
and ( n799 , n120 , n798 ); 
not ( n800 , n120 ); 
not ( n801 , n117 ); 
nand ( n802 , n801 , n73 ); 
and ( n803 , n800 , n802 ); 
or ( n804 , n799 , n803 ); 
not ( n805 , n120 ); 
nand ( n806 , n805 , n41 , n117 ); 
nand ( n807 , n51 , n297 ); 
nand ( n808 , n804 , n806 , n807 ); 
not ( n809 , n808 ); 
not ( n810 , n809 ); 
or ( n811 , n797 , n810 ); 
nand ( n812 , n808 , n321 ); 
nand ( n813 , n811 , n812 ); 
not ( n814 , n813 ); 
not ( n815 , n814 ); 
or ( n816 , n793 , n815 ); 
not ( n817 , n792 ); 
nand ( n818 , n813 , n817 ); 
nand ( n819 , n816 , n818 ); 
not ( n820 , n244 ); 
not ( n821 , n300 ); 
or ( n822 , n820 , n821 ); 
nand ( n823 , n299 , n307 ); 
nand ( n824 , n822 , n823 ); 
not ( n825 , n824 ); 
and ( n826 , n819 , n825 ); 
not ( n827 , n819 ); 
and ( n828 , n827 , n824 ); 
nor ( n829 , n826 , n828 ); 
not ( n830 , n829 ); 
not ( n831 , n830 ); 
or ( n832 , n785 , n831 ); 
and ( n833 , n783 , n829 ); 
nor ( n834 , n833 , n29 ); 
nand ( n835 , n832 , n834 ); 
nand ( n836 , n676 , n768 , n835 ); 
nor ( n837 , n630 , n836 ); 
not ( n838 , n837 ); 
not ( n839 , n23 ); 
or ( n840 , n839 , n747 ); 
nand ( n841 , n21 , n839 ); 
nand ( n842 , n840 , n841 ); 
or ( n843 , n140 , n842 ); 
and ( n844 , n839 , n25 ); 
not ( n845 , n839 ); 
and ( n846 , n845 , n737 ); 
nor ( n847 , n844 , n846 ); 
or ( n848 , n633 , n847 ); 
nand ( n849 , n843 , n848 , n9 ); 
not ( n850 , n849 ); 
not ( n851 , n23 ); 
not ( n852 , n703 ); 
or ( n853 , n851 , n852 ); 
nand ( n854 , n27 , n839 ); 
nand ( n855 , n853 , n854 ); 
not ( n856 , n855 ); 
or ( n857 , n641 , n856 ); 
not ( n858 , n688 ); 
or ( n859 , n839 , n858 ); 
or ( n860 , n22 , n23 ); 
nand ( n861 , n857 , n859 , n860 ); 
not ( n862 , n140 ); 
not ( n863 , n842 ); 
or ( n864 , n862 , n863 ); 
not ( n865 , n141 ); 
and ( n866 , n23 , n476 ); 
not ( n867 , n23 ); 
and ( n868 , n867 , n26 ); 
nor ( n869 , n866 , n868 ); 
nand ( n870 , n865 , n869 ); 
nand ( n871 , n864 , n870 ); 
nor ( n872 , n861 , n871 ); 
not ( n873 , n12 ); 
not ( n874 , n796 ); 
or ( n875 , n873 , n874 ); 
not ( n876 , n12 ); 
nand ( n877 , n13 , n876 ); 
nand ( n878 , n875 , n877 ); 
xnor ( n879 , n878 , n125 ); 
or ( n880 , n142 , n855 ); 
or ( n881 , n865 , n869 ); 
nand ( n882 , n880 , n881 ); 
nor ( n883 , n879 , n882 ); 
and ( n884 , n872 , n883 ); 
and ( n885 , n839 , n24 ); 
not ( n886 , n839 ); 
and ( n887 , n886 , n564 ); 
nor ( n888 , n885 , n887 ); 
nand ( n889 , n322 , n888 ); 
not ( n890 , n322 ); 
not ( n891 , n888 ); 
and ( n892 , n890 , n891 ); 
and ( n893 , n23 , n544 ); 
not ( n894 , n23 ); 
and ( n895 , n894 , n20 ); 
nor ( n896 , n893 , n895 ); 
and ( n897 , n525 , n896 ); 
nor ( n898 , n892 , n897 ); 
not ( n899 , n525 ); 
not ( n900 , n896 ); 
and ( n901 , n899 , n900 ); 
and ( n902 , n633 , n847 ); 
nor ( n903 , n901 , n902 ); 
and ( n904 , n889 , n898 , n903 ); 
nand ( n905 , n850 , n884 , n904 ); 
not ( n906 , n12 ); 
not ( n907 , n424 ); 
or ( n908 , n906 , n907 ); 
nand ( n909 , n15 , n876 ); 
nand ( n910 , n908 , n909 ); 
xnor ( n911 , n910 , n130 ); 
not ( n912 , n12 ); 
not ( n913 , n378 ); 
or ( n914 , n912 , n913 ); 
nand ( n915 , n5 , n876 ); 
nand ( n916 , n914 , n915 ); 
xnor ( n917 , n916 , n129 ); 
nor ( n918 , n911 , n917 ); 
not ( n919 , n12 ); 
not ( n920 , n301 ); 
or ( n921 , n919 , n920 ); 
nand ( n922 , n4 , n876 ); 
nand ( n923 , n921 , n922 ); 
and ( n924 , n923 , n126 ); 
not ( n925 , n923 ); 
and ( n926 , n925 , n653 ); 
nor ( n927 , n924 , n926 ); 
and ( n928 , n12 , n244 ); 
not ( n929 , n12 ); 
and ( n930 , n929 , n14 ); 
nor ( n931 , n928 , n930 ); 
and ( n932 , n931 , n611 ); 
not ( n933 , n931 ); 
and ( n934 , n933 , n128 ); 
nor ( n935 , n932 , n934 ); 
and ( n936 , n918 , n927 , n935 ); 
and ( n937 , n12 , n346 ); 
not ( n938 , n12 ); 
and ( n939 , n938 , n17 ); 
nor ( n940 , n937 , n939 ); 
and ( n941 , n940 , n132 ); 
not ( n942 , n940 ); 
and ( n943 , n942 , n333 ); 
nor ( n944 , n941 , n943 ); 
and ( n945 , n12 , n400 ); 
not ( n946 , n12 ); 
and ( n947 , n946 , n16 ); 
nor ( n948 , n945 , n947 ); 
xor ( n949 , n948 , n131 ); 
nor ( n950 , n944 , n949 ); 
not ( n951 , n23 ); 
not ( n952 , n521 ); 
or ( n953 , n951 , n952 ); 
nand ( n954 , n19 , n839 ); 
nand ( n955 , n953 , n954 ); 
not ( n956 , n955 ); 
or ( n957 , n500 , n956 ); 
or ( n958 , n135 , n955 ); 
not ( n959 , n12 ); 
not ( n960 , n494 ); 
or ( n961 , n959 , n960 ); 
nand ( n962 , n18 , n876 ); 
nand ( n963 , n961 , n962 ); 
nand ( n964 , n134 , n963 ); 
nand ( n965 , n957 , n958 , n964 ); 
and ( n966 , n12 , n448 ); 
and ( n967 , n6 , n876 ); 
nor ( n968 , n966 , n967 ); 
or ( n969 , n432 , n968 ); 
not ( n970 , n963 ); 
nand ( n971 , n473 , n970 ); 
nand ( n972 , n432 , n968 ); 
nand ( n973 , n969 , n971 , n972 ); 
nor ( n974 , n965 , n973 ); 
nand ( n975 , n936 , n950 , n974 ); 
nor ( n976 , n905 , n975 ); 
not ( n977 , n976 ); 
not ( n978 , n808 ); 
or ( n979 , n123 , n978 ); 
not ( n980 , n783 ); 
not ( n981 , n118 ); 
nand ( n982 , n981 , n300 ); 
not ( n983 , n982 ); 
not ( n984 , n825 ); 
or ( n985 , n983 , n984 ); 
not ( n986 , n982 ); 
nand ( n987 , n986 , n824 ); 
nand ( n988 , n985 , n987 ); 
and ( n989 , n988 , n814 ); 
not ( n990 , n988 ); 
and ( n991 , n990 , n813 ); 
nor ( n992 , n989 , n991 ); 
not ( n993 , n992 ); 
not ( n994 , n993 ); 
or ( n995 , n980 , n994 ); 
and ( n996 , n784 , n992 ); 
not ( n997 , n123 ); 
nor ( n998 , n996 , n997 ); 
nand ( n999 , n995 , n998 ); 
nand ( n1000 , n979 , n999 ); 
not ( n1001 , n768 ); 
not ( n1002 , n835 ); 
not ( n1003 , n122 ); 
or ( n1004 , n1003 , n978 ); 
and ( n1005 , n300 , n796 ); 
not ( n1006 , n300 ); 
and ( n1007 , n1006 , n321 ); 
nor ( n1008 , n1005 , n1007 ); 
and ( n1009 , n1008 , n982 ); 
not ( n1010 , n1008 ); 
and ( n1011 , n1010 , n986 ); 
or ( n1012 , n1009 , n1011 ); 
or ( n1013 , n978 , n1012 ); 
and ( n1014 , n978 , n1012 ); 
nor ( n1015 , n1014 , n122 ); 
nand ( n1016 , n1013 , n1015 ); 
nand ( n1017 , n1004 , n1016 ); 
nand ( n1018 , n144 , 1'b1 ); 
xor ( n1019 , n858 , n143 ); 
nand ( n1020 , 1'b1 , n1018 , n1019 ); 
or ( n1021 , n122 , n986 ); 
or ( n1022 , n1003 , n302 ); 
nand ( n1023 , n1021 , n1022 ); 
or ( n1024 , n997 , n986 ); 
or ( n1025 , n123 , n321 ); 
nand ( n1026 , n1024 , n1025 ); 
or ( n1027 , n123 , n302 ); 
or ( n1028 , n997 , n373 ); 
nand ( n1029 , n1027 , n1028 ); 
or ( n1030 , n123 , n307 ); 
not ( n1031 , n424 ); 
or ( n1032 , n997 , n1031 ); 
nand ( n1033 , n1030 , n1032 ); 
not ( n1034 , n1031 ); 
nand ( n1035 , n122 , n321 ); 
nand ( n1036 , n116 , n121 , n28 , n593 ); 
not ( n1037 , n703 ); 
nand ( n1038 , n1 , n3 ); 
nand ( n1039 , n121 , n1038 , n116 , n593 ); 
nor ( n1040 , n591 , n589 ); 
not ( n1041 , n1040 ); 
nand ( n1042 , n7 , n121 ); 
not ( n1043 , n1042 ); 
nand ( n1044 , n1043 , n119 ); 
not ( n1045 , n1042 ); 
nand ( n1046 , n1045 , n147 ); 
not ( n1047 , n542 ); 
nand ( n1048 , n121 , n2 , n11 ); 
nand ( n1049 , n139 , n140 , n141 , n142 ); 
not ( n1050 , n539 ); 
not ( n1051 , n535 ); 
and ( n1052 , n74 , n115 ); 
not ( n1053 , n106 ); 
not ( n1054 , n86 ); 
not ( n1055 , n76 ); 
not ( n1056 , n32 ); 
not ( n1057 , n96 ); 
not ( n1058 , n43 ); 
not ( n1059 , n53 ); 
not ( n1060 , n64 ); 
patch p0 (.t_0(t_0), .g1(n322), .g2(n321), .g3(n435), .g4(n125));
endmodule 

