module patch (t_0, t_1, t_2, t_3, t_4, t_5, t_6, t_7, t_8, t_9, t_10, t_11, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18;
output t_0, t_1, t_2, t_3, t_4, t_5, t_6, t_7, t_8, t_9, t_10, t_11;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882;

nor ( w8882 , w1407 , w1395 );
and ( w1 , w8792 , g2 );
and ( w2 , w1 , w8735 );
and ( w3 , w2 , w8860 );
and ( w4 , w3 , w8769 );
and ( w5 , w4 , w8845 );
nor ( w6 , w5 , g5 );
nor ( w7 , w6 , g7 );
nor ( w8 , w7 , g4 );
not ( w9 , w8 );
and ( w10 , w9 , g8 );
nor ( w11 , w10 , g7 );
and ( w12 , w11 , g8 );
and ( w13 , w8735 , g8 );
and ( w14 , w8769 , w13 );
and ( w15 , w8742 , g8 );
and ( w16 , w5546 , g8 );
nor ( w17 , g5 , g9 );
not ( w18 , w16 );
and ( w19 , w18 , w17 );
nor ( w20 , w19 , g5 );
not ( w21 , w20 );
and ( w22 , w14 , w21 );
not ( w23 , w22 );
and ( w24 , w23 , g8 );
and ( w25 , w24 , w8742 );
and ( w26 , w25 , w8769 );
nor ( w27 , g4 , g3 );
not ( w28 , w26 );
and ( w29 , w28 , w27 );
nor ( w30 , w29 , g4 );
nor ( w31 , w12 , w30 );
and ( w32 , w31 , g10 );
and ( w33 , g10 , w8792 );
and ( w34 , w32 , w33 );
not ( w35 , w34 );
and ( w36 , w35 , g10 );
nor ( w37 , w36 , g6 );
and ( w38 , w37 , w8765 );
and ( w39 , w38 , g2 );
nor ( w40 , g1 , g2 );
and ( w41 , w40 , w8765 );
and ( w42 , w41 , w8845 );
and ( w43 , w42 , w8860 );
and ( w44 , w43 , w8735 );
and ( w45 , w44 , w8742 );
and ( w46 , w45 , g10 );
and ( w47 , w46 , w8769 );
nor ( w48 , w47 , g5 );
nor ( w49 , w48 , g7 );
and ( w50 , w49 , g10 );
nor ( w51 , w50 , g7 );
nor ( w52 , w51 , g6 );
and ( w53 , w52 , w13 );
not ( w54 , w53 );
and ( w55 , w54 , g8 );
and ( w56 , w8837 , g8 );
not ( w57 , w56 );
and ( w58 , w57 , g8 );
nor ( w59 , g5 , g7 );
and ( w60 , w58 , w59 );
nor ( w61 , w60 , g7 );
and ( w62 , w61 , w59 );
not ( w63 , w62 );
and ( w64 , w63 , g12 );
and ( w65 , w64 , w8742 );
not ( w66 , w65 );
and ( w67 , w66 , w17 );
nor ( w68 , w67 , g5 );
nor ( w69 , w68 , g3 );
nor ( w70 , g5 , w59 );
and ( w71 , w70 , w8742 );
not ( w72 , w71 );
and ( w73 , w72 , g10 );
and ( w74 , w73 , g8 );
not ( w75 , w74 );
and ( w76 , w75 , g8 );
and ( w77 , w17 , w8742 );
nor ( w78 , w77 , g5 );
and ( w79 , w78 , w8742 );
not ( w80 , w79 );
and ( w81 , w80 , g8 );
not ( w82 , w81 );
and ( w83 , w82 , g8 );
nor ( w84 , w76 , w83 );
and ( w85 , w84 , w8735 );
and ( w86 , w85 , w7783 );
and ( w87 , w86 , w8860 );
and ( w88 , w87 , g10 );
and ( w89 , w88 , w8765 );
and ( w90 , w89 , w8792 );
and ( w91 , w69 , w90 );
nor ( w92 , g3 , g10 );
nor ( w93 , w91 , w92 );
nor ( w94 , w93 , g9 );
and ( w95 , w94 , w7783 );
and ( w96 , w95 , w8819 );
and ( w97 , w96 , g14 );
and ( w98 , w97 , w8792 );
not ( w99 , w55 );
and ( w100 , w99 , w98 );
and ( w101 , w100 , g10 );
nor ( w102 , w101 , w92 );
nor ( w103 , w102 , g6 );
nor ( w104 , g6 , g2 );
and ( w105 , w103 , w104 );
and ( w106 , w105 , w8765 );
and ( w107 , w106 , w8819 );
and ( w108 , w107 , g14 );
and ( w109 , w108 , w8792 );
nor ( w110 , g4 , w109 );
not ( w111 , w92 );
and ( w112 , w110 , w111 );
nor ( w113 , w112 , g6 );
and ( w114 , w113 , w8765 );
and ( w115 , w114 , w7783 );
and ( w116 , w115 , w8819 );
and ( w117 , w116 , g14 );
and ( w118 , w117 , g15 );
and ( w119 , w8728 , g14 );
and ( w120 , w119 , g15 );
and ( w121 , w8735 , g10 );
nor ( w122 , g1 , g15 );
and ( w123 , w8735 , w122 );
and ( w124 , w123 , w8742 );
and ( w125 , w124 , g11 );
and ( w126 , w125 , g2 );
nor ( w127 , w121 , w126 );
and ( w128 , g5 , g3 );
not ( w129 , w128 );
and ( w130 , w127 , w129 );
nor ( w131 , w130 , g14 );
and ( w132 , w8769 , g3 );
not ( w133 , w132 );
and ( w134 , w133 , w122 );
and ( w135 , w134 , g14 );
and ( w136 , w135 , w8828 );
nor ( w137 , w131 , w136 );
nor ( w138 , w137 , g12 );
and ( w139 , w138 , w8860 );
and ( w140 , w139 , w8828 );
and ( w141 , w140 , w8819 );
and ( w142 , w141 , g6 );
and ( w143 , w142 , g11 );
and ( w144 , w143 , g2 );
and ( w145 , w144 , w8792 );
nor ( w146 , w120 , w145 );
nor ( w147 , w146 , g16 );
and ( w148 , w147 , w8819 );
and ( w149 , w148 , g6 );
and ( w150 , g3 , w8828 );
and ( w151 , w150 , w8819 );
and ( w152 , w151 , w8742 );
and ( w153 , w152 , w8765 );
and ( w154 , w153 , w8728 );
and ( w155 , w154 , w8845 );
and ( w156 , w155 , g2 );
and ( w157 , w156 , g11 );
and ( w158 , w157 , w8792 );
nor ( w159 , w149 , w158 );
not ( w160 , w159 );
and ( w161 , w160 , g11 );
and ( w162 , g11 , w8819 );
and ( w163 , w162 , w8828 );
and ( w164 , w123 , w8845 );
and ( w165 , w164 , g12 );
and ( w166 , w165 , w8860 );
and ( w167 , w166 , w8837 );
and ( w168 , w167 , w8819 );
and ( w169 , w168 , w7783 );
and ( w170 , w169 , w8765 );
and ( w171 , w170 , w8828 );
nor ( w172 , g4 , w171 );
nor ( w173 , w172 , g11 );
and ( w174 , w173 , w8819 );
and ( w175 , w174 , w7783 );
and ( w176 , w175 , w8765 );
and ( w177 , w176 , w8828 );
and ( w178 , w177 , w8792 );
nor ( w179 , w163 , w178 );
not ( w180 , w179 );
and ( w181 , w180 , g4 );
not ( w182 , w123 );
and ( w183 , w182 , g14 );
nor ( w184 , w183 , g3 );
and ( w185 , w184 , w8819 );
and ( w186 , w185 , w8828 );
and ( w187 , w186 , w7783 );
and ( w188 , w187 , w8860 );
and ( w189 , w188 , w8765 );
and ( w190 , w189 , w8792 );
and ( w191 , w190 , g12 );
and ( w192 , w191 , w7141 );
and ( w193 , w192 , w8845 );
and ( w194 , w193 , w8837 );
and ( w195 , w190 , w8845 );
and ( w196 , w195 , g11 );
nor ( w197 , w196 , w178 );
not ( w198 , w194 );
and ( w199 , w198 , w197 );
not ( w200 , w181 );
and ( w201 , w200 , w199 );
nor ( w202 , w201 , g2 );
and ( w203 , w202 , w8765 );
and ( w204 , w203 , w8792 );
nor ( w205 , w161 , w204 );
not ( w206 , w205 );
and ( w207 , w206 , g2 );
nor ( w208 , w207 , w204 );
not ( w209 , w118 );
and ( w210 , w209 , w208 );
nor ( w211 , w210 , g16 );
nor ( w212 , w39 , w211 );
and ( w213 , g14 , w8168 );
and ( w214 , w212 , w213 );
not ( w215 , w121 );
and ( w216 , w215 , g10 );
not ( w217 , w216 );
and ( w218 , w217 , g15 );
and ( w219 , w218 , w8860 );
and ( w220 , w184 , w8860 );
and ( w221 , w220 , w8792 );
and ( w222 , w219 , w221 );
nor ( w223 , w222 , w123 );
and ( w224 , w8730 , g15 );
and ( w225 , w224 , g7 );
and ( w226 , w225 , w8769 );
nor ( w227 , w223 , w226 );
and ( w228 , w227 , g11 );
and ( w229 , w228 , w8860 );
and ( w230 , w229 , w8819 );
not ( w231 , w230 );
and ( w232 , w231 , g11 );
and ( w233 , w232 , w8728 );
not ( w234 , w233 );
and ( w235 , w234 , w221 );
and ( w236 , w235 , w8845 );
and ( w237 , w236 , g2 );
not ( w238 , w237 );
and ( w239 , w238 , w208 );
nor ( w240 , g1 , g6 );
and ( w241 , w240 , g2 );
and ( w242 , w241 , w8765 );
and ( w243 , w242 , w8860 );
and ( w244 , w243 , w8735 );
and ( w245 , w244 , g10 );
and ( w246 , w245 , w59 );
nor ( w247 , w246 , g5 );
and ( w248 , w247 , w8860 );
and ( w249 , w248 , w8742 );
nor ( w250 , w249 , g6 );
and ( w251 , w250 , g2 );
and ( w252 , g11 , w251 );
and ( w253 , w252 , w8769 );
nor ( w254 , w253 , g5 );
nor ( w255 , w254 , g7 );
nor ( w256 , w255 , g4 );
not ( w257 , w256 );
and ( w258 , w257 , g8 );
nor ( w259 , w258 , g7 );
not ( w260 , w259 );
and ( w261 , w260 , g8 );
not ( w262 , w261 );
and ( w263 , w262 , g8 );
and ( w264 , w121 , w59 );
nor ( w265 , w264 , g5 );
nor ( w266 , w265 , g4 );
and ( w267 , w266 , w8765 );
and ( w268 , w267 , w8735 );
and ( w269 , w268 , w8845 );
and ( w270 , w8735 , g7 );
nor ( w271 , w269 , w270 );
nor ( w272 , w271 , g6 );
nor ( w273 , g4 , w272 );
nor ( w274 , w273 , g6 );
not ( w275 , w263 );
and ( w276 , w275 , w274 );
and ( w277 , w276 , g10 );
and ( w278 , w277 , w33 );
nor ( w279 , w278 , w92 );
nor ( w280 , w279 , g6 );
and ( w281 , w280 , w8765 );
and ( w282 , w281 , g2 );
and ( w283 , w282 , w8819 );
and ( w284 , w283 , g15 );
nor ( w285 , w284 , w211 );
not ( w286 , w285 );
and ( w287 , w286 , g14 );
and ( w288 , w287 , g15 );
and ( w289 , w1 , w8765 );
and ( w290 , w289 , w8860 );
and ( w291 , w290 , w8735 );
and ( w292 , w291 , w8837 );
nor ( w293 , w292 , w230 );
not ( w294 , w293 );
and ( w295 , w294 , g2 );
and ( w296 , w295 , w8728 );
and ( w297 , w8735 , g4 );
and ( w298 , w297 , w122 );
and ( w299 , g5 , g7 );
and ( w300 , w299 , w8730 );
not ( w301 , w300 );
and ( w302 , w301 , w2 );
and ( w303 , w302 , w7141 );
and ( w304 , w303 , g15 );
nor ( w305 , w298 , w304 );
not ( w306 , w305 );
and ( w307 , w306 , g4 );
nor ( w308 , w307 , w221 );
nor ( w309 , w308 , g6 );
not ( w310 , w309 );
and ( w311 , w310 , w208 );
not ( w312 , w311 );
and ( w313 , w312 , g2 );
and ( w314 , w313 , g11 );
nor ( w315 , w123 , w297 );
nor ( w316 , w315 , g6 );
and ( w317 , w316 , g2 );
and ( w318 , w317 , w8837 );
and ( w319 , w318 , g12 );
and ( w320 , w319 , w8819 );
and ( w321 , w320 , w8792 );
nor ( w322 , w314 , w321 );
not ( w323 , w322 );
and ( w324 , w323 , g12 );
and ( w325 , w324 , w8819 );
and ( w326 , w325 , w7997 );
and ( w327 , w326 , w8828 );
not ( w328 , w327 );
and ( w329 , w328 , w208 );
and ( w330 , w8728 , g4 );
and ( w331 , w1037 , w329 );
nor ( w332 , w331 , g6 );
not ( w333 , w332 );
and ( w334 , w333 , w208 );
not ( w335 , w334 );
and ( w336 , w335 , g2 );
and ( w337 , w336 , w8735 );
and ( w338 , w337 , w8765 );
and ( w339 , w338 , w8819 );
and ( w340 , w339 , w7997 );
and ( w341 , w340 , w8828 );
and ( w342 , w341 , w8792 );
not ( w343 , w342 );
and ( w344 , w329 , w343 );
not ( w345 , w344 );
and ( w346 , w345 , g2 );
and ( w347 , w346 , w8735 );
and ( w348 , w347 , w8765 );
not ( w349 , w348 );
and ( w350 , w349 , w208 );
nor ( w351 , w350 , w213 );
nor ( w352 , w296 , w351 );
not ( w353 , w352 );
and ( w354 , w353 , w27 );
nor ( w355 , w354 , w342 );
nor ( w356 , w355 , g6 );
not ( w357 , w356 );
and ( w358 , w357 , w208 );
not ( w359 , w358 );
and ( w360 , w359 , g2 );
nor ( w361 , g3 , g9 );
and ( w362 , w360 , w361 );
not ( w363 , w362 );
and ( w364 , w363 , w208 );
nor ( w365 , w364 , g13 );
and ( w366 , w365 , w7997 );
and ( w367 , w366 , w8828 );
nor ( w368 , w288 , w367 );
nor ( w369 , w368 , g16 );
not ( w370 , w369 );
and ( w371 , w239 , w370 );
not ( w372 , w371 );
and ( w373 , w372 , w361 );
not ( w374 , w373 );
and ( w375 , w374 , w208 );
nor ( w376 , w369 , g12 );
and ( w377 , w376 , w8837 );
and ( w378 , w8765 , w377 );
nor ( w379 , w375 , w378 );
and ( w380 , w379 , w27 );
and ( w381 , g14 , g15 );
nor ( w382 , w380 , w381 );
nor ( w383 , w382 , g3 );
and ( w384 , w383 , w8819 );
nor ( w385 , w384 , w369 );
nor ( w386 , w385 , g16 );
nor ( w387 , w386 , w381 );
nor ( w388 , w214 , w387 );
nor ( w389 , w247 , g7 );
nor ( w390 , w389 , g4 );
not ( w391 , w390 );
and ( w392 , w391 , g8 );
nor ( w393 , w392 , g7 );
not ( w394 , w393 );
and ( w395 , w394 , w13 );
not ( w396 , w395 );
and ( w397 , w396 , g8 );
not ( w398 , w397 );
and ( w399 , w398 , w274 );
and ( w400 , w8845 , g2 );
and ( w401 , w399 , w400 );
nor ( w402 , w401 , w211 );
not ( w403 , w402 );
and ( w404 , w403 , g10 );
not ( w405 , w404 );
and ( w406 , w405 , w213 );
and ( w407 , w221 , w8845 );
nor ( w408 , g1 , g9 );
and ( w409 , w407 , w408 );
and ( w410 , w409 , w436 );
nor ( w411 , w410 , w342 );
not ( w412 , w411 );
and ( w413 , w412 , g2 );
nor ( w414 , w413 , w369 );
and ( w415 , w414 , w7934 );
not ( w416 , w415 );
and ( w417 , w416 , g10 );
and ( w418 , w92 , w8765 );
and ( w419 , w418 , g2 );
nor ( w420 , w419 , w211 );
and ( w421 , w420 , w213 );
and ( w422 , w230 , w8845 );
not ( w423 , w422 );
and ( w424 , w423 , g11 );
and ( w425 , w424 , w8728 );
and ( w426 , w418 , w8819 );
and ( w427 , w426 , w8860 );
and ( w428 , w427 , w8828 );
not ( w429 , w428 );
and ( w430 , w429 , g12 );
nor ( w431 , w430 , g10 );
and ( w432 , w431 , w8735 );
and ( w433 , w432 , w8828 );
not ( w434 , w425 );
and ( w435 , w434 , w433 );
not ( w436 , w377 );
and ( w437 , w435 , w436 );
not ( w438 , w437 );
and ( w439 , w438 , w208 );
not ( w440 , w439 );
and ( w441 , w440 , w361 );
and ( w442 , w441 , w408 );
and ( w443 , w442 , w27 );
nor ( w444 , w443 , w381 );
nor ( w445 , w444 , g10 );
and ( w446 , w445 , w8735 );
and ( w447 , w446 , w8819 );
nor ( w448 , w447 , w369 );
nor ( w449 , w448 , g16 );
nor ( w450 , w449 , w381 );
nor ( w451 , w421 , w450 );
and ( w452 , w451 , w8730 );
and ( w453 , w452 , w8735 );
and ( w454 , w453 , w8819 );
nor ( w455 , w454 , w369 );
nor ( w456 , w455 , g16 );
nor ( w457 , w417 , w456 );
nor ( w458 , w457 , g3 );
and ( w459 , w458 , w8819 );
nor ( w460 , w459 , w369 );
nor ( w461 , w460 , g16 );
not ( w462 , w406 );
and ( w463 , w462 , w461 );
and ( w464 , w463 , w33 );
nor ( w465 , w464 , w456 );
not ( w466 , w465 );
nand ( t_0 , w388 , w466 );
and ( w467 , g4 , w8845 );
and ( w468 , w467 , w8765 );
and ( w469 , w468 , g15 );
and ( w470 , w469 , w8819 );
and ( w471 , w408 , w8845 );
and ( w472 , w471 , w8860 );
and ( w473 , w472 , w8742 );
and ( w474 , w473 , g8 );
and ( w475 , w474 , w8769 );
and ( w476 , w8845 , g5 );
and ( w477 , w476 , w8735 );
nor ( w478 , w475 , w477 );
not ( w479 , w478 );
and ( w480 , w479 , w27 );
nor ( w481 , w480 , g4 );
not ( w482 , w481 );
and ( w483 , w482 , g10 );
and ( w484 , w483 , w33 );
and ( w485 , w484 , w13 );
nor ( w486 , w485 , w270 );
and ( w487 , w92 , w8828 );
and ( w488 , w486 , w972 );
nor ( w489 , g3 , g8 );
and ( w490 , w488 , w970 );
not ( w491 , w490 );
and ( w492 , w491 , w400 );
and ( w493 , w492 , w8765 );
and ( w494 , w493 , w8819 );
and ( w495 , w187 , w8792 );
and ( w496 , w495 , g12 );
and ( w497 , w496 , g15 );
and ( w498 , w497 , w8845 );
and ( w499 , w498 , w8837 );
and ( w500 , g15 , w8735 );
and ( w501 , w500 , w8845 );
and ( w502 , w501 , w8837 );
and ( w503 , w502 , g16 );
and ( w504 , w503 , w8819 );
and ( w505 , w504 , w8765 );
and ( w506 , w505 , w7783 );
and ( w507 , w506 , w7997 );
and ( w508 , w476 , g3 );
and ( w509 , w508 , g11 );
and ( w510 , w509 , w8765 );
and ( w511 , w510 , w8792 );
nor ( w512 , g1 , g3 );
and ( w513 , w512 , g6 );
and ( w514 , w513 , w7783 );
and ( w515 , w514 , w8765 );
and ( w516 , w515 , w8860 );
nor ( w517 , w511 , w516 );
and ( w518 , w408 , w8860 );
and ( w519 , w518 , w7783 );
and ( w520 , w519 , g3 );
and ( w521 , w520 , w122 );
not ( w522 , w521 );
and ( w523 , w522 , g14 );
not ( w524 , w523 );
and ( w525 , w524 , w520 );
and ( w526 , g6 , g3 );
and ( w527 , w525 , w526 );
not ( w528 , w527 );
and ( w529 , w517 , w528 );
nor ( w530 , w529 , g12 );
nor ( w531 , w530 , w178 );
not ( w532 , w531 );
and ( w533 , w532 , g11 );
nor ( w534 , w533 , w178 );
nor ( w535 , w534 , g13 );
and ( w536 , w535 , w7783 );
and ( w537 , w536 , w8828 );
and ( w538 , w495 , w8845 );
and ( w539 , w538 , g11 );
nor ( w540 , w539 , w178 );
nor ( w541 , w540 , g9 );
and ( w542 , w541 , w7997 );
nor ( w543 , w537 , w542 );
not ( w544 , w507 );
and ( w545 , w544 , w543 );
nor ( w546 , w545 , w213 );
nor ( w547 , w499 , w546 );
and ( w548 , w547 , w545 );
nor ( w549 , w548 , g9 );
and ( w550 , w549 , w7997 );
nor ( w551 , g4 , g12 );
and ( w552 , w291 , w8728 );
not ( w553 , w552 );
and ( w554 , w551 , w553 );
nor ( w555 , w554 , g13 );
and ( w556 , w555 , w8735 );
and ( w557 , w556 , w8845 );
and ( w558 , w557 , w8792 );
and ( w559 , w558 , g2 );
and ( w560 , w559 , w8828 );
nor ( w561 , g3 , g12 );
nor ( w562 , w561 , w270 );
and ( w563 , w562 , w967 );
and ( w564 , w563 , w970 );
and ( w565 , w46 , g8 );
and ( w566 , w565 , w8769 );
and ( w567 , w566 , g12 );
not ( w568 , w567 );
and ( w569 , w564 , w568 );
nor ( w570 , w569 , g6 );
nor ( w571 , g4 , w567 );
nor ( w572 , w571 , g6 );
nor ( w573 , w572 , w487 );
nor ( w574 , w573 , g9 );
and ( w575 , w574 , g15 );
and ( w576 , w575 , w7783 );
and ( w577 , w576 , w8828 );
nor ( w578 , w570 , w577 );
and ( w579 , w578 , w972 );
nor ( w580 , w579 , g9 );
and ( w581 , w580 , w8819 );
and ( w582 , w581 , g15 );
and ( w583 , w582 , g14 );
and ( w584 , w583 , w7783 );
and ( w585 , w584 , w8828 );
nor ( w586 , w585 , w549 );
nor ( w587 , w586 , g11 );
nor ( w588 , w587 , w549 );
not ( w589 , w560 );
and ( w590 , w589 , w588 );
nor ( w591 , w590 , w213 );
not ( w592 , w591 );
and ( w593 , w592 , w588 );
nor ( w594 , w593 , g11 );
nor ( w595 , w550 , w594 );
and ( w596 , w595 , w588 );
not ( w597 , w494 );
and ( w598 , w597 , w596 );
not ( w599 , w598 );
and ( w600 , w599 , g14 );
and ( w601 , w600 , g15 );
not ( w602 , w601 );
and ( w603 , w602 , w596 );
nor ( w604 , w603 , g11 );
and ( w605 , w604 , w8828 );
and ( w606 , w330 , w8845 );
and ( w607 , w606 , w7997 );
and ( w608 , w607 , w8819 );
and ( w609 , w608 , w8792 );
and ( w610 , w609 , w8828 );
and ( w611 , w610 , w8730 );
and ( w612 , g5 , w967 );
not ( w613 , w612 );
and ( w614 , w613 , g10 );
and ( w615 , w614 , w8845 );
and ( w616 , w615 , w8735 );
nor ( w617 , w611 , w616 );
nor ( w618 , w617 , g13 );
and ( w619 , w618 , w8735 );
and ( w620 , w619 , w7997 );
and ( w621 , w620 , w8765 );
and ( w622 , w621 , w8828 );
nor ( w623 , w622 , w610 );
not ( w624 , w623 );
and ( w625 , w624 , g11 );
and ( w626 , w625 , w8728 );
nor ( w627 , w527 , w549 );
nor ( w628 , w627 , g16 );
nor ( w629 , g2 , w628 );
nor ( w630 , w629 , g12 );
and ( w631 , w630 , g6 );
and ( w632 , w8728 , g2 );
nor ( w633 , w632 , w550 );
nor ( w634 , w633 , g6 );
and ( w635 , w634 , w8819 );
and ( w636 , w635 , g11 );
and ( w637 , w636 , w7997 );
and ( w638 , w637 , w8765 );
nor ( w639 , w631 , w638 );
not ( w640 , w639 );
and ( w641 , w640 , g3 );
and ( w642 , w641 , g11 );
nor ( w643 , g12 , w527 );
and ( w644 , w643 , g3 );
and ( w645 , w644 , w7783 );
and ( w646 , w645 , w8860 );
and ( w647 , w646 , w8769 );
and ( w648 , w647 , w8819 );
and ( w649 , w648 , g6 );
not ( w650 , w649 );
and ( w651 , w650 , g11 );
and ( w652 , w651 , w8828 );
and ( w653 , w642 , w652 );
not ( w654 , w605 );
and ( w655 , w654 , w588 );
and ( w656 , w655 , w8730 );
and ( w657 , w656 , g15 );
and ( w658 , w657 , w8860 );
and ( w659 , w658 , w8742 );
and ( w660 , g15 , w8860 );
nor ( w661 , w660 , w122 );
nor ( w662 , w661 , g7 );
nor ( w663 , w662 , g7 );
and ( w664 , w663 , w8860 );
nor ( w665 , w659 , w664 );
and ( w666 , w665 , g6 );
and ( w667 , w666 , w8728 );
and ( w668 , w655 , w1037 );
not ( w669 , w622 );
and ( w670 , w668 , w669 );
nor ( w671 , w670 , g10 );
nor ( w672 , w671 , w616 );
nor ( w673 , w672 , g6 );
and ( w674 , w673 , w8819 );
not ( w675 , w674 );
and ( w676 , w675 , w655 );
nor ( w677 , w676 , g3 );
and ( w678 , w677 , g11 );
and ( w679 , w678 , w652 );
nor ( w680 , w679 , w550 );
nor ( w681 , w680 , w213 );
and ( w682 , w681 , w8765 );
and ( w683 , w682 , w8828 );
not ( w684 , w683 );
and ( w685 , w655 , w684 );
not ( w686 , w667 );
and ( w687 , w686 , w685 );
not ( w688 , w687 );
and ( w689 , w688 , g2 );
and ( w690 , g2 , w8735 );
and ( w691 , w689 , w690 );
nor ( w692 , w691 , w550 );
not ( w693 , w692 );
and ( w694 , w693 , g6 );
nor ( w695 , w694 , w683 );
nor ( w696 , w695 , g13 );
not ( w697 , w696 );
and ( w698 , w697 , w655 );
nor ( w699 , w698 , g3 );
and ( w700 , w699 , w361 );
and ( w701 , w700 , g11 );
and ( w702 , w701 , w652 );
nor ( w703 , w702 , w550 );
nor ( w704 , w703 , w213 );
and ( w705 , w704 , w8828 );
nor ( w706 , w653 , w705 );
not ( w707 , w550 );
and ( w708 , w706 , w707 );
nor ( w709 , w708 , g13 );
not ( w710 , w709 );
and ( w711 , w710 , w655 );
nor ( w712 , w711 , w213 );
and ( w713 , w712 , w8792 );
and ( w714 , w713 , w8765 );
and ( w715 , w714 , w8828 );
nor ( w716 , w549 , w715 );
and ( w717 , w716 , w655 );
not ( w718 , w626 );
and ( w719 , w718 , w717 );
not ( w720 , w719 );
and ( w721 , w720 , g2 );
not ( w722 , w721 );
and ( w723 , w722 , w717 );
nor ( w724 , w723 , g3 );
nor ( w725 , w724 , w715 );
and ( w726 , w725 , w655 );
nor ( w727 , w726 , w213 );
and ( w728 , w727 , w8765 );
and ( w729 , w728 , w8828 );
nor ( w730 , w605 , w729 );
and ( w731 , w730 , w717 );
and ( w732 , w244 , w8769 );
and ( w733 , w732 , g8 );
and ( w734 , w733 , g10 );
and ( w735 , w734 , w8742 );
and ( w736 , w735 , g14 );
and ( w737 , w736 , g15 );
and ( w738 , w737 , g12 );
and ( w739 , w738 , w8819 );
not ( w740 , w739 );
and ( w741 , w740 , w655 );
not ( w742 , w741 );
and ( w743 , w742 , g11 );
not ( w744 , w743 );
and ( w745 , w744 , w655 );
nor ( w746 , w745 , g16 );
not ( w747 , w746 );
and ( w748 , w747 , w655 );
and ( w749 , w731 , w748 );
and ( w750 , g12 , w655 );
not ( w751 , w750 );
and ( w752 , w751 , g3 );
and ( w753 , w752 , w8845 );
and ( w754 , w753 , g15 );
and ( w755 , w754 , g2 );
nor ( w756 , g3 , w516 );
nor ( w757 , w756 , g12 );
nor ( w758 , w487 , g12 );
and ( w759 , w16 , w8742 );
not ( w760 , w759 );
and ( w761 , w760 , w33 );
and ( w762 , w761 , w17 );
not ( w763 , w762 );
and ( w764 , w763 , g10 );
and ( w765 , w764 , w8769 );
and ( w766 , w1847 , g5 );
nor ( w767 , w766 , g10 );
nor ( w768 , w767 , g10 );
and ( w769 , w768 , g7 );
nor ( w770 , w769 , g3 );
and ( w771 , w770 , w7783 );
and ( w772 , w771 , w8860 );
and ( w773 , w5412 , w772 );
and ( w774 , w773 , w8792 );
not ( w775 , w758 );
and ( w776 , w775 , w774 );
nor ( w777 , w776 , g4 );
nor ( w778 , w777 , g2 );
and ( w779 , w8860 , g10 );
and ( w780 , w779 , g12 );
and ( w781 , w780 , w7783 );
and ( w782 , w59 , g8 );
and ( w783 , w781 , w782 );
not ( w784 , w783 );
and ( w785 , w778 , w784 );
and ( w786 , w785 , w8735 );
and ( w787 , w786 , g6 );
not ( w788 , w782 );
and ( w789 , w270 , w788 );
and ( w790 , w789 , w8728 );
and ( w791 , w616 , g7 );
not ( w792 , w791 );
and ( w793 , w792 , g7 );
not ( w794 , w793 );
and ( w795 , w794 , w17 );
and ( w796 , w616 , g5 );
nor ( w797 , w795 , w796 );
nor ( w798 , w797 , g3 );
and ( w799 , w798 , w8860 );
and ( w800 , w799 , w8845 );
and ( w801 , w800 , g8 );
and ( w802 , w616 , w8767 );
nor ( w803 , w801 , w802 );
nor ( w804 , w803 , w782 );
and ( w805 , w804 , w33 );
and ( w806 , w487 , w8860 );
nor ( w807 , w805 , w806 );
and ( w808 , w738 , w8828 );
not ( w809 , w808 );
and ( w810 , w807 , w809 );
not ( w811 , w810 );
and ( w812 , w811 , w27 );
and ( w813 , w812 , g12 );
and ( w814 , w813 , w8845 );
and ( w815 , w814 , g14 );
and ( w816 , w815 , g15 );
and ( w817 , w816 , w8819 );
and ( w818 , w817 , w8828 );
nor ( w819 , w790 , w818 );
and ( w820 , w819 , w8860 );
nor ( w821 , w820 , g6 );
and ( w822 , w821 , g14 );
and ( w823 , w822 , g15 );
and ( w824 , w823 , w8819 );
and ( w825 , w824 , w8828 );
nor ( w826 , w787 , w825 );
not ( w827 , w826 );
and ( w828 , w827 , g14 );
and ( w829 , w828 , g15 );
and ( w830 , w829 , w8819 );
and ( w831 , w830 , w8828 );
not ( w832 , w831 );
and ( w833 , w832 , w655 );
not ( w834 , w833 );
and ( w835 , w834 , g11 );
not ( w836 , w835 );
and ( w837 , w836 , w655 );
and ( w838 , w8728 , g3 );
and ( w839 , w838 , w7783 );
and ( w840 , w839 , g11 );
not ( w841 , w840 );
and ( w842 , w841 , w655 );
nor ( w843 , w842 , g13 );
not ( w844 , w843 );
and ( w845 , w844 , w731 );
nor ( w846 , w845 , g9 );
and ( w847 , w846 , g14 );
not ( w848 , w847 );
and ( w849 , w848 , w731 );
nor ( w850 , w849 , g16 );
not ( w851 , w850 );
and ( w852 , w837 , w851 );
and ( w853 , w852 , w8860 );
nor ( w854 , w853 , g6 );
and ( w855 , w854 , g15 );
and ( w856 , w855 , w7783 );
and ( w857 , w856 , g11 );
not ( w858 , w857 );
and ( w859 , w858 , w655 );
nor ( w860 , w859 , g13 );
not ( w861 , w860 );
and ( w862 , w861 , w731 );
nor ( w863 , w862 , g9 );
and ( w864 , w863 , g14 );
not ( w865 , w864 );
and ( w866 , w865 , w731 );
nor ( w867 , w866 , g16 );
not ( w868 , w867 );
and ( w869 , w868 , w655 );
and ( w870 , w869 , w837 );
and ( w871 , w757 , w8730 );
and ( w872 , w871 , w7783 );
and ( w873 , w872 , w8765 );
not ( w874 , w873 );
and ( w875 , w870 , w874 );
not ( w876 , w875 );
and ( w877 , w876 , g6 );
nor ( w878 , w877 , w867 );
not ( w879 , w878 );
and ( w880 , w879 , g15 );
and ( w881 , w880 , w7783 );
and ( w882 , w881 , g11 );
not ( w883 , w882 );
and ( w884 , w883 , w655 );
nor ( w885 , w884 , g13 );
not ( w886 , w885 );
and ( w887 , w886 , w731 );
nor ( w888 , w887 , g9 );
and ( w889 , w888 , g14 );
not ( w890 , w889 );
and ( w891 , w890 , w731 );
nor ( w892 , w891 , g16 );
nor ( w893 , w757 , w892 );
not ( w894 , w893 );
and ( w895 , w894 , g6 );
nor ( w896 , w895 , w867 );
not ( w897 , w896 );
and ( w898 , w897 , g15 );
and ( w899 , w898 , w7783 );
and ( w900 , w899 , g11 );
not ( w901 , w900 );
and ( w902 , w901 , w655 );
nor ( w903 , w902 , g13 );
not ( w904 , w903 );
and ( w905 , w904 , w731 );
nor ( w906 , w905 , g9 );
and ( w907 , w906 , g14 );
not ( w908 , w907 );
and ( w909 , w908 , w731 );
nor ( w910 , w909 , g16 );
not ( w911 , w910 );
and ( w912 , w911 , w655 );
not ( w913 , w755 );
and ( w914 , w913 , w912 );
not ( w915 , w914 );
and ( w916 , w915 , g11 );
not ( w917 , w916 );
and ( w918 , w917 , w655 );
nor ( w919 , w918 , g13 );
and ( w920 , w919 , w8765 );
and ( w921 , w920 , g14 );
not ( w922 , w921 );
and ( w923 , w922 , w731 );
nor ( w924 , w923 , g16 );
not ( w925 , w924 );
and ( w926 , w655 , w925 );
and ( w927 , g12 , w926 );
not ( w928 , w927 );
and ( w929 , w928 , g6 );
nor ( w930 , w929 , w924 );
not ( w931 , w930 );
and ( w932 , w931 , g15 );
and ( w933 , w932 , g2 );
not ( w934 , w933 );
and ( w935 , w934 , w912 );
not ( w936 , w935 );
and ( w937 , w936 , g11 );
not ( w938 , w937 );
and ( w939 , w938 , w655 );
nor ( w940 , w939 , g13 );
and ( w941 , w940 , w8765 );
and ( w942 , w941 , g14 );
not ( w943 , w942 );
and ( w944 , w943 , w731 );
nor ( w945 , w944 , g16 );
not ( w946 , w945 );
and ( w947 , w946 , w912 );
and ( w948 , w749 , w947 );
not ( w949 , w470 );
and ( w950 , w949 , w948 );
not ( w951 , w950 );
and ( w952 , w951 , g14 );
not ( w953 , w952 );
and ( w954 , w953 , w731 );
nor ( w955 , w954 , g16 );
and ( w956 , w955 , w8845 );
and ( w957 , w956 , g15 );
not ( w958 , w957 );
and ( w959 , w958 , w948 );
not ( w960 , w959 );
and ( w961 , w960 , g11 );
not ( w962 , w961 );
and ( w963 , w962 , w655 );
and ( w964 , w963 , w8860 );
not ( w965 , w964 );
and ( w966 , w965 , g11 );
not ( w967 , w477 );
and ( w968 , g12 , w967 );
and ( w969 , w968 , w5920 );
not ( w970 , w489 );
and ( w971 , w969 , w970 );
not ( w972 , w487 );
and ( w973 , w971 , w972 );
not ( w974 , w973 );
and ( w975 , w974 , g2 );
and ( w976 , w975 , w8845 );
nor ( w977 , w976 , w585 );
nor ( w978 , w977 , g11 );
not ( w979 , w978 );
and ( w980 , w979 , w963 );
nor ( w981 , w980 , g6 );
and ( w982 , w981 , g14 );
and ( w983 , w982 , g15 );
and ( w984 , w617 , g11 );
not ( w985 , w984 );
and ( w986 , w985 , w560 );
not ( w987 , w986 );
and ( w988 , w987 , w963 );
nor ( w989 , w988 , w213 );
not ( w990 , w989 );
and ( w991 , w990 , w963 );
nor ( w992 , w616 , w487 );
nor ( w993 , w992 , g12 );
nor ( w994 , w993 , w818 );
not ( w995 , w818 );
and ( w996 , w995 , w963 );
and ( w997 , w994 , w996 );
and ( w998 , w997 , w8860 );
nor ( w999 , w998 , g6 );
and ( w1000 , w999 , g14 );
and ( w1001 , w1000 , w8765 );
and ( w1002 , w1001 , w8819 );
not ( w1003 , w1002 );
and ( w1004 , w1003 , w963 );
nor ( w1005 , w1004 , g16 );
and ( w1006 , w1005 , w8728 );
nor ( w1007 , w1006 , w818 );
not ( w1008 , w1007 );
and ( w1009 , w1008 , g11 );
nor ( w1010 , w1009 , g4 );
nor ( w1011 , w1010 , g6 );
not ( w1012 , w1011 );
and ( w1013 , w1012 , w963 );
not ( w1014 , w1013 );
and ( w1015 , w1014 , g14 );
and ( w1016 , w1015 , g15 );
and ( w1017 , w487 , w8742 );
and ( w1018 , w806 , g5 );
and ( w1019 , w487 , w122 );
nor ( w1020 , w1018 , w1019 );
nor ( w1021 , w1020 , g4 );
and ( w1022 , w1021 , w8728 );
and ( w1023 , w1019 , g12 );
and ( w1024 , w477 , w8742 );
and ( w1025 , w487 , w8769 );
nor ( w1026 , w1024 , w1025 );
not ( w1027 , w806 );
and ( w1028 , w1026 , w1027 );
not ( w1029 , w1028 );
and ( w1030 , w1029 , g12 );
and ( w1031 , w1030 , w8730 );
and ( w1032 , w1031 , w8845 );
and ( w1033 , w1032 , g2 );
and ( w1034 , w1033 , w8792 );
and ( w1035 , w1034 , w8828 );
nor ( w1036 , w1023 , w1035 );
not ( w1037 , w330 );
and ( w1038 , w1036 , w1037 );
nor ( w1039 , w1038 , g10 );
and ( w1040 , w1039 , w8845 );
and ( w1041 , w1040 , g2 );
and ( w1042 , w1041 , w7997 );
and ( w1043 , w1042 , w8819 );
and ( w1044 , w1043 , w8792 );
and ( w1045 , w1044 , w8828 );
nor ( w1046 , w1022 , w1045 );
not ( w1047 , w616 );
and ( w1048 , w1046 , w1047 );
nor ( w1049 , w1048 , g6 );
and ( w1050 , w1049 , w8735 );
and ( w1051 , w1050 , g2 );
and ( w1052 , w1051 , w7997 );
and ( w1053 , w1052 , w8819 );
and ( w1054 , w1053 , w8792 );
and ( w1055 , w1054 , w8828 );
nor ( w1056 , w1017 , w1055 );
not ( w1057 , w1019 );
and ( w1058 , w1056 , w1057 );
nor ( w1059 , w1058 , g4 );
and ( w1060 , w1059 , w8728 );
nor ( w1061 , w1060 , w1045 );
nor ( w1062 , w1061 , g10 );
nor ( w1063 , w1062 , w616 );
and ( w1064 , w1063 , g11 );
not ( w1065 , w1064 );
and ( w1066 , w1065 , w560 );
not ( w1067 , w1066 );
and ( w1068 , w1067 , w963 );
nor ( w1069 , w1068 , g6 );
and ( w1070 , w1069 , w7997 );
and ( w1071 , w1070 , g2 );
nor ( w1072 , w487 , w831 );
not ( w1073 , w1072 );
and ( w1074 , w1073 , g14 );
and ( w1075 , w1074 , g15 );
and ( w1076 , w1075 , w8765 );
and ( w1077 , w1076 , w8819 );
not ( w1078 , w1077 );
and ( w1079 , w1078 , w963 );
nor ( w1080 , w1079 , g16 );
nor ( w1081 , w1080 , w1005 );
not ( w1082 , w1081 );
and ( w1083 , w1082 , g11 );
and ( w1084 , w1083 , g14 );
and ( w1085 , w1084 , g15 );
not ( w1086 , w1085 );
and ( w1087 , w1086 , w963 );
nor ( w1088 , w1087 , g2 );
not ( w1089 , w1088 );
and ( w1090 , w1089 , w963 );
nor ( w1091 , w1090 , g16 );
nor ( w1092 , w1071 , w1091 );
nor ( w1093 , w1092 , g9 );
not ( w1094 , w1093 );
and ( w1095 , w1094 , w963 );
not ( w1096 , w1016 );
and ( w1097 , w1096 , w1095 );
not ( w1098 , w1097 );
and ( w1099 , w1098 , g2 );
nor ( w1100 , w1099 , w1091 );
nor ( w1101 , w1100 , g9 );
and ( w1102 , w1101 , w8819 );
not ( w1103 , w1102 );
and ( w1104 , w1103 , w963 );
nor ( w1105 , w1104 , g16 );
not ( w1106 , w1105 );
and ( w1107 , w991 , w1106 );
nor ( w1108 , w1107 , g9 );
not ( w1109 , w1108 );
and ( w1110 , w1109 , w963 );
not ( w1111 , w983 );
and ( w1112 , w1111 , w1110 );
nor ( w1113 , w1112 , g9 );
and ( w1114 , w1113 , w8819 );
not ( w1115 , w1114 );
and ( w1116 , w1115 , w963 );
nor ( w1117 , w1116 , g16 );
nor ( w1118 , w966 , w1117 );
nor ( w1119 , w1118 , g6 );
and ( w1120 , w1119 , g14 );
and ( w1121 , w1120 , g15 );
not ( w1122 , w1121 );
and ( w1123 , w1122 , w1110 );
nor ( w1124 , w1123 , g9 );
and ( w1125 , w1124 , w8819 );
not ( w1126 , w1125 );
and ( w1127 , w1126 , w963 );
nor ( w1128 , w1127 , g1 );
and ( w1129 , w1128 , w8828 );
not ( w1130 , w1129 );
and ( w1131 , w1130 , w1110 );
and ( w1132 , w8828 , w1131 );
and ( w1133 , w1276 , g15 );
not ( w1134 , w1133 );
and ( w1135 , w1134 , w1131 );
nor ( w1136 , w1135 , w213 );
and ( w1137 , w1136 , w8735 );
and ( w1138 , w1137 , w8837 );
not ( w1139 , w1138 );
and ( w1140 , w1131 , w1139 );
nor ( w1141 , w1140 , g6 );
and ( w1142 , w1141 , g12 );
not ( w1143 , w1142 );
and ( w1144 , w1143 , w1131 );
not ( w1145 , w1144 );
and ( w1146 , w1145 , g2 );
and ( w1147 , w1146 , w8837 );
not ( w1148 , w1147 );
and ( w1149 , w1148 , w1131 );
nor ( w1150 , w1149 , g9 );
not ( w1151 , w1150 );
and ( w1152 , w1131 , w1151 );
and ( w1153 , w1131 , w8728 );
nor ( w1154 , w1153 , w1132 );
and ( w1155 , w1154 , w8730 );
and ( w1156 , w1155 , w8735 );
and ( w1157 , w1156 , g2 );
not ( w1158 , w1157 );
and ( w1159 , w1158 , w1131 );
nor ( w1160 , w1159 , g11 );
not ( w1161 , w1160 );
and ( w1162 , w1161 , w1131 );
and ( w1163 , w1152 , w1162 );
nor ( w1164 , w1163 , g9 );
and ( w1165 , w1164 , w8735 );
and ( w1166 , w1165 , g2 );
and ( w1167 , w1166 , w8837 );
not ( w1168 , w1167 );
and ( w1169 , w1131 , w1168 );
and ( w1170 , w1276 , w477 );
and ( w1171 , w1170 , w8819 );
not ( w1172 , w1171 );
and ( w1173 , w1131 , w1172 );
not ( w1174 , w1173 );
and ( w1175 , w1174 , g14 );
and ( w1176 , w1175 , g15 );
not ( w1177 , w1176 );
and ( w1178 , w1177 , w1131 );
nor ( w1179 , w1178 , g11 );
not ( w1180 , w1179 );
and ( w1181 , w1180 , w1131 );
and ( w1182 , w1131 , g11 );
nor ( w1183 , w1132 , g1 );
and ( w1184 , w1183 , w8735 );
and ( w1185 , w1184 , w8767 );
and ( w1186 , w1185 , w8845 );
nor ( w1187 , w1132 , g3 );
and ( w1188 , w1187 , w8730 );
and ( w1189 , w1188 , w8767 );
and ( w1190 , w1186 , w1189 );
and ( w1191 , w1190 , g2 );
and ( w1192 , w1191 , g14 );
and ( w1193 , w1192 , g15 );
not ( w1194 , w1193 );
and ( w1195 , w1194 , w1131 );
nor ( w1196 , w1195 , g5 );
and ( w1197 , w1196 , w8742 );
not ( w1198 , w1197 );
and ( w1199 , w1198 , g12 );
not ( w1200 , w1199 );
and ( w1201 , w1200 , w59 );
and ( w1202 , w1201 , w8730 );
and ( w1203 , w1202 , w1276 );
and ( w1204 , w1203 , g2 );
and ( w1205 , w1204 , w8845 );
and ( w1206 , w1205 , w8765 );
and ( w1207 , w1206 , w27 );
and ( w1208 , w1207 , w408 );
not ( w1209 , w1208 );
and ( w1210 , w1131 , w1209 );
not ( w1211 , w1210 );
and ( w1212 , w1211 , g12 );
not ( w1213 , w1212 );
and ( w1214 , w1213 , w1131 );
not ( w1215 , w1214 );
and ( w1216 , w1215 , g2 );
and ( w1217 , w1216 , w8765 );
nor ( w1218 , w1217 , g11 );
and ( w1219 , w1218 , w1131 );
nor ( w1220 , g9 , g8 );
nor ( w1221 , w1220 , g8 );
not ( w1222 , w1221 );
and ( w1223 , w1222 , w59 );
and ( w1224 , w1223 , w8860 );
nor ( w1225 , w1224 , g7 );
and ( w1226 , w1225 , w8769 );
nor ( w1227 , w1226 , w1132 );
and ( w1228 , w1227 , w8735 );
nor ( w1229 , w1228 , g4 );
nor ( w1230 , w1229 , w1132 );
nor ( w1231 , w1221 , w1132 );
and ( w1232 , w1231 , w8765 );
and ( w1233 , w1230 , w1232 );
and ( w1234 , g10 , w8767 );
nor ( w1235 , w1234 , g8 );
and ( w1236 , w6486 , w27 );
and ( w1237 , w1236 , w8845 );
nor ( w1238 , w1237 , g4 );
not ( w1239 , w1238 );
and ( w1240 , w1233 , w1239 );
and ( w1241 , w1240 , w33 );
nor ( w1242 , w1241 , w1188 );
and ( w1243 , w104 , w8767 );
nor ( w1244 , g7 , g4 );
and ( w1245 , w1243 , w1244 );
nor ( w1246 , w1245 , g8 );
and ( w1247 , w1246 , w8860 );
and ( w1248 , g10 , w8769 );
not ( w1249 , w1247 );
and ( w1250 , w1249 , w1248 );
not ( w1251 , w1250 );
and ( w1252 , w1251 , g10 );
nor ( w1253 , w1252 , g9 );
nor ( w1254 , w1253 , g5 );
and ( w1255 , w1254 , w8742 );
nor ( w1256 , w1255 , g3 );
and ( w1257 , w1256 , w1276 );
not ( w1258 , w1242 );
and ( w1259 , w1258 , w1257 );
nor ( w1260 , g2 , g3 );
and ( w1261 , w1259 , w1260 );
and ( w1262 , w1261 , w8845 );
and ( w1263 , w1262 , w408 );
and ( w1264 , g12 , w8742 );
and ( w1265 , w1264 , w8860 );
and ( w1266 , w1265 , g10 );
and ( w1267 , w1266 , w8769 );
and ( w1268 , w1267 , w8767 );
nor ( w1269 , w1268 , g6 );
and ( w1270 , w1263 , w1269 );
and ( w1271 , w1270 , g11 );
and ( w1272 , w1271 , g13 );
not ( w1273 , w1272 );
and ( w1274 , w1131 , w1273 );
and ( w1275 , w1276 , g4 );
not ( w1276 , w1132 );
and ( w1277 , w40 , w1276 );
and ( w1278 , w1277 , w8765 );
and ( w1279 , w1278 , w8767 );
and ( w1280 , w1279 , w8860 );
and ( w1281 , w1280 , w8845 );
and ( w1282 , w1281 , w59 );
and ( w1283 , w1282 , w8730 );
nor ( w1284 , w1283 , g7 );
and ( w1285 , w1284 , w8767 );
and ( w1286 , w1285 , w8769 );
nor ( w1287 , w1286 , w1132 );
and ( w1288 , w1287 , w8730 );
and ( w1289 , w1288 , w7783 );
and ( w1290 , w1289 , w104 );
and ( w1291 , w1290 , w8765 );
and ( w1292 , w1187 , w1291 );
and ( w1293 , w1292 , w8860 );
and ( w1294 , w1293 , w408 );
nor ( w1295 , w1275 , w1294 );
nor ( w1296 , w1295 , g10 );
and ( w1297 , w1296 , w7783 );
and ( w1298 , w1297 , w8845 );
and ( w1299 , w1298 , w8765 );
and ( w1300 , w1187 , w1299 );
not ( w1301 , w1300 );
and ( w1302 , w1301 , w1131 );
not ( w1303 , w1302 );
and ( w1304 , w1303 , g14 );
and ( w1305 , w1304 , g15 );
and ( w1306 , w1305 , w7783 );
and ( w1307 , w1306 , w8845 );
not ( w1308 , w1307 );
and ( w1309 , w1131 , w1308 );
nor ( w1310 , w1309 , g11 );
not ( w1311 , w1310 );
and ( w1312 , w1311 , w1131 );
not ( w1313 , w1312 );
and ( w1314 , w1313 , g13 );
not ( w1315 , w1314 );
and ( w1316 , w1315 , w1131 );
and ( w1317 , w1274 , w1316 );
not ( w1318 , w1317 );
and ( w1319 , w1318 , g14 );
and ( w1320 , w1319 , g15 );
not ( w1321 , w1320 );
and ( w1322 , w1321 , w1131 );
and ( w1323 , w1219 , w1322 );
not ( w1324 , w1323 );
and ( w1325 , w1324 , g13 );
not ( w1326 , w1325 );
and ( w1327 , w1326 , w1131 );
nor ( w1328 , w1182 , w1327 );
not ( w1329 , w1328 );
and ( w1330 , w1329 , w1322 );
and ( w1331 , w1181 , w1330 );
nor ( w1332 , w1331 , g9 );
not ( w1333 , w1332 );
and ( w1334 , w1333 , w1131 );
nor ( w1335 , w1334 , g2 );
not ( w1336 , w1335 );
and ( w1337 , w1336 , w1131 );
nor ( w1338 , w1337 , g11 );
not ( w1339 , w1338 );
and ( w1340 , w1339 , w1131 );
and ( w1341 , w1340 , w1330 );
nor ( w1342 , w1341 , g9 );
not ( w1343 , w1342 );
and ( w1344 , w1169 , w1343 );
nor ( w1345 , w1344 , g13 );
not ( w1346 , w1345 );
and ( t_1 , w1346 , w1330 );
and ( w1347 , w241 , g10 );
and ( w1348 , g8 , g9 );
not ( w1349 , w1348 );
and ( w1350 , w1349 , g8 );
not ( w1351 , w1350 );
and ( w1352 , w1351 , w241 );
and ( w1353 , w1 , w8730 );
and ( w1354 , w1353 , g8 );
not ( w1355 , w1354 );
and ( w1356 , w1355 , g8 );
not ( w1357 , w1356 );
and ( w1358 , w1357 , w241 );
and ( w1359 , w1352 , w1358 );
and ( w1360 , w1359 , w8730 );
and ( w1361 , w8730 , g9 );
and ( w1362 , w1360 , w1361 );
nor ( w1363 , w1347 , w1362 );
not ( w1364 , w1363 );
and ( w1365 , w1364 , g9 );
and ( w1366 , g17 , w8767 );
and ( w1367 , w1366 , w8730 );
not ( w1368 , w1367 );
and ( w1369 , w1368 , w241 );
and ( w1370 , w1369 , w8765 );
not ( w1371 , w1370 );
and ( w1372 , w1371 , g14 );
and ( w1373 , w1372 , w8168 );
and ( w1374 , w1373 , g13 );
nor ( w1375 , w1374 , g6 );
and ( w1376 , w1375 , g2 );
and ( w1377 , w1376 , w8792 );
nor ( w1378 , w1377 , g16 );
not ( w1379 , w1365 );
and ( w1380 , w1379 , w1378 );
nor ( w1381 , w1380 , g6 );
not ( w1382 , w1381 );
and ( w1383 , w1382 , g11 );
nor ( w1384 , w381 , g9 );
and ( w1385 , w1384 , w8735 );
and ( w1386 , w1385 , w8728 );
and ( w1387 , w1386 , g4 );
and ( w1388 , w1387 , w8769 );
and ( w1389 , w1388 , w8742 );
and ( w1390 , w1389 , g13 );
and ( w1391 , w1390 , w7783 );
and ( w1392 , w1391 , w8845 );
and ( w1393 , w1392 , w8837 );
and ( w1394 , w1393 , g16 );
and ( w1395 , w1394 , w8792 );
nor ( w1396 , w1383 , w1395 );
not ( w1397 , w1396 );
and ( w1398 , w1397 , g13 );
not ( w1399 , w1398 );
and ( w1400 , w1399 , w400 );
nor ( w1401 , w1400 , g6 );
not ( w1402 , w1401 );
and ( w1403 , w1402 , g2 );
not ( w1404 , w1403 );
and ( w1405 , w1404 , g2 );
nor ( w1406 , w1405 , g1 );
nor ( w1407 , w1406 , g1 );
or ( t_2 , w1407 , w1395 );
nor ( w1408 , w1361 , g10 );
not ( w1409 , w1408 );
and ( w1410 , w1409 , g2 );
and ( w1411 , w1410 , w8845 );
nor ( w1412 , w1411 , g6 );
and ( w1413 , w1412 , g13 );
nor ( w1414 , g10 , g8 );
and ( w1415 , w1414 , g16 );
and ( w1416 , w1415 , g2 );
and ( w1417 , w1416 , w8845 );
and ( w1418 , w1417 , w8837 );
and ( w1419 , w1418 , w8792 );
and ( w1420 , w1419 , g9 );
and ( w1421 , w27 , g12 );
and ( w1422 , w1421 , w8742 );
and ( w1423 , w1422 , w8769 );
nor ( w1424 , w1423 , g10 );
and ( w1425 , w1424 , w8767 );
and ( w1426 , w1425 , g13 );
nor ( w1427 , w1244 , g7 );
and ( w1428 , w1427 , w8860 );
nor ( w1429 , w1428 , g9 );
nor ( w1430 , w1429 , g1 );
and ( w1431 , w1430 , g6 );
and ( w1432 , w1431 , w8837 );
and ( w1433 , w1432 , g16 );
nor ( w1434 , w1426 , w1433 );
not ( w1435 , w1434 );
and ( w1436 , w1435 , g14 );
nor ( w1437 , w1436 , w1433 );
not ( w1438 , w1437 );
and ( w1439 , w1438 , g16 );
and ( w1440 , w1439 , w8765 );
and ( w1441 , w1440 , g2 );
nor ( w1442 , w1441 , w1433 );
nor ( w1443 , w1442 , g6 );
nor ( w1444 , w1443 , w1433 );
nor ( w1445 , w1444 , g11 );
and ( w1446 , w1445 , w8792 );
nor ( w1447 , w1420 , w1446 );
not ( w1448 , w1413 );
and ( w1449 , w1448 , w1447 );
not ( w1450 , w1449 );
and ( w1451 , w1450 , g2 );
and ( w1452 , w1451 , g11 );
and ( w1453 , w1452 , g16 );
and ( w1454 , w1453 , g14 );
and ( w1455 , w1454 , w8168 );
not ( w1456 , w1455 );
and ( w1457 , w1456 , w1447 );
nor ( w1458 , w1457 , g1 );
and ( w1459 , w8765 , g13 );
nor ( w1460 , w1459 , g10 );
nor ( w1461 , w1460 , g10 );
not ( w1462 , w1461 );
and ( w1463 , w1462 , g6 );
not ( w1464 , w1463 );
and ( w1465 , w1464 , g6 );
and ( w1466 , w1465 , w7783 );
and ( w1467 , w1466 , g11 );
and ( w1468 , w1467 , g16 );
and ( w1469 , w1468 , g14 );
and ( w1470 , w1469 , w8168 );
and ( w1471 , w1470 , w8792 );
nor ( w1472 , w1458 , w1471 );
nor ( w1473 , g1 , g8 );
and ( w1474 , w1473 , w1423 );
and ( w1475 , w1474 , w8730 );
nor ( w1476 , w1475 , g8 );
nor ( w1477 , w1476 , g10 );
and ( w1478 , w1477 , w408 );
and ( w1479 , w1478 , w7783 );
nor ( w1480 , w1479 , g2 );
nor ( w1481 , w1480 , g10 );
nor ( w1482 , w1481 , g11 );
and ( w1483 , w1482 , g16 );
and ( w1484 , w1483 , g14 );
and ( w1485 , w1484 , w8168 );
nor ( w1486 , w1485 , g1 );
and ( w1487 , w1486 , w8765 );
and ( w1488 , w1487 , g12 );
and ( w1489 , g6 , w7783 );
and ( w1490 , w1488 , w1489 );
nor ( w1491 , w1490 , g2 );
nor ( w1492 , w1491 , g10 );
nor ( w1493 , w1492 , g10 );
not ( w1494 , w1493 );
and ( w1495 , w1494 , g6 );
not ( w1496 , w1495 );
and ( w1497 , w1496 , g6 );
and ( w1498 , w1497 , w8837 );
and ( w1499 , w1498 , g16 );
and ( w1500 , w1499 , g14 );
and ( w1501 , w1500 , w8168 );
nor ( w1502 , w1501 , w1433 );
and ( w1503 , w1502 , w8792 );
and ( w1504 , w1503 , w8730 );
nor ( w1505 , w1504 , g10 );
not ( w1506 , w1505 );
and ( w1507 , w1506 , g6 );
not ( w1508 , w1507 );
and ( w1509 , w1508 , g6 );
not ( w1510 , w1509 );
and ( w1511 , w1510 , w1447 );
nor ( w1512 , w1511 , g1 );
not ( w1513 , w1512 );
nand ( t_3 , w1472 , w1513 );
and ( w1514 , w1 , g3 );
and ( w1515 , w8845 , g10 );
and ( w1516 , w8792 , g6 );
and ( w1517 , w1516 , g2 );
and ( w1518 , g9 , w1414 );
nor ( w1519 , w1518 , g8 );
and ( w1520 , w6151 , w1519 );
nor ( w1521 , w1520 , g1 );
and ( w1522 , w4929 , g14 );
and ( w1523 , w1522 , w8168 );
nor ( w1524 , w1523 , g1 );
not ( w1525 , w1524 );
and ( w1526 , w1525 , g11 );
and ( w1527 , w8882 , g10 );
nor ( w1528 , w1527 , g11 );
nor ( w1529 , w1526 , w1528 );
and ( w1530 , w1529 , w400 );
and ( w1531 , w40 , w4939 );
nor ( w1532 , w1530 , w1531 );
nor ( w1533 , w1532 , g1 );
not ( w1534 , w1533 );
and ( w1535 , w1534 , g16 );
and ( w1536 , w471 , w8735 );
and ( w1537 , w1536 , g5 );
nor ( w1538 , w1537 , w17 );
and ( w1539 , w1536 , g7 );
not ( w1540 , w1539 );
and ( w1541 , w1540 , g7 );
not ( w1542 , w1541 );
and ( w1543 , w1542 , g8 );
and ( w1544 , w512 , w8767 );
nor ( w1545 , w1543 , w1544 );
nor ( w1546 , w1545 , g1 );
and ( w1547 , w1546 , w8765 );
and ( w1548 , w1547 , w8845 );
not ( w1549 , w1538 );
and ( w1550 , w1549 , w1548 );
and ( w1551 , w1550 , w33 );
and ( w1552 , w512 , w8730 );
nor ( w1553 , w1551 , w1552 );
nor ( w1554 , w1553 , g9 );
nor ( w1555 , w122 , g6 );
and ( w1556 , w1555 , w8860 );
and ( w1557 , w1556 , w8735 );
and ( w1558 , w1557 , w8765 );
and ( w1559 , w1558 , g2 );
and ( w1560 , w1559 , w8819 );
and ( w1561 , w1560 , w7141 );
and ( w1562 , w1561 , w8730 );
and ( w1563 , w1562 , w8728 );
and ( w1564 , w1563 , w8837 );
and ( w1565 , w1564 , w8792 );
and ( w1566 , w1565 , g16 );
nor ( w1567 , w1395 , w1566 );
and ( w1568 , w1554 , w1567 );
and ( w1569 , w1568 , w8845 );
nor ( w1570 , w1430 , w1569 );
not ( w1571 , w1570 );
and ( w1572 , w1571 , g2 );
not ( w1573 , w1519 );
and ( w1574 , w40 , w1573 );
and ( w1575 , w7783 , g18 );
not ( w1576 , w1575 );
and ( w1577 , w1576 , g18 );
nor ( w1578 , w1577 , g10 );
and ( w1579 , g9 , w8767 );
and ( w1580 , w1578 , w1579 );
nor ( w1581 , w1580 , g10 );
and ( w1582 , w1581 , w8767 );
nor ( w1583 , g6 , w1582 );
and ( w1584 , w1574 , w1583 );
and ( w1585 , w1584 , w8730 );
and ( w1586 , w1585 , g9 );
nor ( w1587 , w770 , g3 );
nor ( w1588 , w1587 , g1 );
nor ( w1589 , w512 , g1 );
nor ( w1590 , w500 , g1 );
not ( w1591 , w1590 );
and ( w1592 , w1591 , w1567 );
and ( w1593 , w1592 , w8765 );
and ( w1594 , w1593 , w8735 );
and ( w1595 , w1594 , g10 );
and ( w1596 , w1595 , g7 );
and ( w1597 , w1596 , g2 );
not ( w1598 , w1597 );
and ( w1599 , w1598 , g11 );
nor ( w1600 , w1599 , g4 );
and ( w1601 , w1600 , g2 );
and ( w1602 , w1601 , w8735 );
nor ( w1603 , g4 , w1602 );
nor ( w1604 , w1603 , g12 );
nor ( w1605 , w122 , w1594 );
nor ( w1606 , w1605 , g9 );
and ( w1607 , w1606 , w8792 );
and ( w1608 , w1607 , w8735 );
nor ( w1609 , g5 , g4 );
nor ( w1610 , w1609 , g5 );
not ( w1611 , w1610 );
and ( w1612 , w1608 , w1611 );
and ( w1613 , w8769 , g7 );
not ( w1614 , w661 );
and ( w1615 , w1614 , w1613 );
nor ( w1616 , w1615 , g5 );
not ( w1617 , w1616 );
and ( w1618 , w1612 , w1617 );
and ( w1619 , g15 , w8769 );
not ( w1620 , w1619 );
and ( w1621 , w1618 , w1620 );
and ( w1622 , w1621 , g7 );
and ( w1623 , w1622 , g2 );
not ( w1624 , w1623 );
and ( w1625 , w1624 , g11 );
nor ( w1626 , w1625 , g4 );
and ( w1627 , w1626 , w361 );
and ( w1628 , w1627 , g2 );
and ( w1629 , w1628 , w8792 );
and ( w1630 , w1629 , g7 );
and ( w1631 , w1630 , w8845 );
nor ( w1632 , g4 , w1631 );
nor ( w1633 , w1632 , g12 );
and ( w1634 , w1594 , g15 );
nor ( w1635 , w1634 , w122 );
nor ( w1636 , w1635 , g3 );
and ( w1637 , w1636 , g4 );
and ( w1638 , w1637 , w408 );
not ( w1639 , w768 );
and ( w1640 , w1639 , w1638 );
and ( w1641 , w1588 , w8168 );
not ( w1642 , w1641 );
and ( w1643 , w1642 , g2 );
nor ( w1644 , w123 , g1 );
not ( w1645 , w1644 );
and ( w1646 , w1645 , w1567 );
and ( w1647 , w1646 , w7783 );
and ( w1648 , w1647 , w8735 );
nor ( w1649 , w1643 , w1648 );
nor ( w1650 , w1649 , g18 );
and ( w1651 , g1 , g2 );
nor ( w1652 , w1651 , g13 );
and ( w1653 , g5 , w8742 );
nor ( w1654 , g7 , w1653 );
nor ( w1655 , w1654 , g15 );
nor ( w1656 , w1655 , g10 );
nor ( w1657 , w1656 , w1654 );
and ( w1658 , w1657 , w7141 );
and ( w1659 , w1655 , g14 );
nor ( w1660 , w1658 , w1659 );
nor ( w1661 , w1660 , w299 );
and ( w1662 , w1661 , w8728 );
and ( w1663 , w1662 , w8765 );
and ( w1664 , w1663 , g3 );
and ( w1665 , w2777 , g12 );
and ( w1666 , w1665 , g7 );
and ( w1667 , w1666 , w7141 );
and ( w1668 , w1667 , g3 );
and ( w1669 , w1421 , w8833 );
and ( w1670 , w1421 , g10 );
and ( w1671 , w1670 , w8735 );
and ( w1672 , w1671 , w8828 );
nor ( w1673 , w1669 , w1672 );
nor ( w1674 , w1673 , g14 );
and ( w1675 , w1674 , w8828 );
nor ( w1676 , w1668 , w1675 );
and ( w1677 , g12 , g7 );
and ( w1678 , w1677 , g3 );
nor ( w1679 , w1678 , w1421 );
nor ( w1680 , w1679 , g4 );
and ( w1681 , w1680 , w8833 );
and ( w1682 , w1681 , g14 );
and ( w1683 , w1682 , w8792 );
and ( w1684 , w1683 , w8828 );
not ( w1685 , w1684 );
and ( w1686 , w1676 , w1685 );
nor ( w1687 , w1686 , g9 );
and ( w1688 , w1687 , w8792 );
and ( w1689 , w1688 , w8828 );
nor ( w1690 , w1664 , w1689 );
not ( w1691 , w1690 );
and ( w1692 , w1691 , g6 );
not ( w1693 , w1692 );
and ( w1694 , w1693 , w1567 );
nor ( w1695 , w1694 , g2 );
and ( w1696 , w1695 , w8792 );
not ( w1697 , w1696 );
and ( w1698 , w1697 , w1567 );
not ( w1699 , w1698 );
and ( w1700 , w1699 , g11 );
and ( w1701 , w1700 , g13 );
and ( w1702 , w1701 , w8828 );
and ( w1703 , w1653 , g12 );
and ( w1704 , w1703 , w8833 );
nor ( w1705 , w1704 , g10 );
not ( w1706 , w1705 );
and ( w1707 , w1706 , w1703 );
and ( w1708 , w1707 , w7141 );
and ( w1709 , w1708 , g11 );
and ( w1710 , w1709 , w8792 );
and ( w1711 , w1710 , w7783 );
and ( w1712 , w1711 , g13 );
and ( w1713 , w1712 , w8828 );
and ( w1714 , w1713 , w8860 );
and ( w1715 , w1714 , g3 );
and ( w1716 , w1715 , w8765 );
not ( w1717 , w1716 );
and ( w1718 , w1717 , w1567 );
and ( w1719 , w59 , g4 );
and ( w1720 , w1719 , w8728 );
and ( w1721 , w1720 , w8735 );
and ( w1722 , w1721 , g11 );
not ( w1723 , w1722 );
and ( w1724 , w1718 , w1723 );
nor ( w1725 , w1724 , g14 );
and ( w1726 , w1703 , w8860 );
and ( w1727 , w1726 , g3 );
and ( w1728 , w1727 , w8765 );
and ( w1729 , w1728 , g11 );
and ( w1730 , w1729 , w8792 );
and ( w1731 , w1730 , g13 );
and ( w1732 , w1731 , w8828 );
and ( w1733 , w1732 , w8833 );
and ( w1734 , w1733 , g14 );
and ( w1735 , w1734 , w7783 );
nor ( w1736 , w1725 , w1735 );
nor ( w1737 , w1736 , g9 );
not ( w1738 , w1737 );
and ( w1739 , w1738 , w1567 );
not ( w1740 , w1739 );
and ( w1741 , w1740 , g6 );
not ( w1742 , w1741 );
and ( w1743 , w1742 , w1567 );
nor ( w1744 , w1743 , g1 );
and ( w1745 , w1744 , w7783 );
and ( w1746 , w1745 , g13 );
and ( w1747 , w1746 , w8828 );
not ( w1748 , w1747 );
and ( w1749 , w1748 , w1567 );
not ( w1750 , w1702 );
and ( w1751 , w1750 , w1749 );
not ( w1752 , w1652 );
and ( w1753 , w1752 , w1751 );
nor ( w1754 , w1753 , g16 );
and ( w1755 , w1588 , w1754 );
and ( w1756 , w1755 , g2 );
and ( w1757 , w8168 , w1567 );
and ( w1758 , w1757 , w1751 );
not ( w1759 , w1756 );
and ( w1760 , w1759 , w1758 );
nor ( w1761 , w1760 , w381 );
not ( w1762 , w1761 );
and ( w1763 , w1762 , g9 );
nor ( w1764 , w1763 , w1594 );
not ( w1765 , w1764 );
and ( w1766 , w1765 , g12 );
and ( w1767 , w1766 , w8845 );
and ( w1768 , w1767 , w8735 );
nor ( w1769 , w1768 , g13 );
not ( w1770 , w1769 );
and ( w1771 , w1770 , w1751 );
nor ( w1772 , w1771 , g16 );
not ( w1773 , w1650 );
and ( w1774 , w1773 , w1772 );
not ( w1775 , w1774 );
and ( w1776 , w1775 , g12 );
and ( w1777 , w1776 , w8845 );
and ( w1778 , w1777 , w8735 );
and ( w1779 , w1778 , w8860 );
and ( w1780 , w1779 , g2 );
and ( w1781 , w1608 , g11 );
nor ( w1782 , w1781 , g4 );
and ( w1783 , w1782 , w8728 );
and ( w1784 , w1594 , w8769 );
nor ( w1785 , w1784 , w1648 );
and ( w1786 , w770 , g5 );
not ( w1787 , w1786 );
and ( w1788 , w1785 , w1787 );
nor ( w1789 , w1788 , g9 );
and ( w1790 , w1789 , w7783 );
not ( w1791 , w1783 );
and ( w1792 , w1791 , w1790 );
nor ( w1793 , w1792 , w381 );
nor ( w1794 , w1793 , g1 );
and ( w1795 , w1794 , w8735 );
nor ( w1796 , w1780 , w1795 );
nor ( w1797 , w381 , g1 );
not ( w1798 , w1797 );
and ( w1799 , w1798 , w1567 );
and ( w1800 , w1799 , w7783 );
and ( w1801 , w1800 , w8845 );
nor ( w1802 , w381 , w1801 );
nor ( w1803 , w1802 , g1 );
nor ( w1804 , w1803 , w381 );
and ( w1805 , w838 , w8860 );
and ( w1806 , w1805 , w8769 );
and ( w1807 , w1806 , w8742 );
and ( w1808 , w1807 , g6 );
and ( w1809 , w1808 , w8765 );
nor ( w1810 , w381 , w1809 );
nor ( w1811 , w1810 , g1 );
and ( w1812 , w1811 , w8735 );
nor ( w1813 , w1801 , w1812 );
and ( w1814 , g11 , w7141 );
and ( w1815 , w1814 , g15 );
and ( w1816 , w1815 , w8730 );
and ( w1817 , w1816 , g4 );
and ( w1818 , w1817 , w299 );
and ( w1819 , w1818 , g12 );
nor ( w1820 , g14 , g12 );
and ( w1821 , w1820 , g15 );
and ( w1822 , w1821 , w8730 );
and ( w1823 , w1822 , w8860 );
and ( w1824 , w1823 , w8769 );
nor ( w1825 , w1819 , w1824 );
not ( w1826 , w1825 );
and ( w1827 , w1826 , g2 );
and ( w1828 , w1827 , w1567 );
and ( w1829 , w1828 , w8845 );
and ( w1830 , w1813 , w1948 );
nor ( w1831 , w1830 , g9 );
and ( w1832 , w1831 , w8792 );
nor ( w1833 , w1832 , w381 );
not ( w1834 , w1833 );
and ( w1835 , w1834 , g7 );
and ( w1836 , w1835 , w8735 );
not ( w1837 , w1836 );
and ( w1838 , w1804 , w1837 );
and ( w1839 , w1796 , w1838 );
nor ( w1840 , w1839 , g1 );
nor ( w1841 , w1840 , g1 );
nor ( w1842 , w1841 , g3 );
and ( w1843 , w1842 , g7 );
nor ( w1844 , g4 , g2 );
nor ( w1845 , w1844 , g4 );
and ( w1846 , g4 , g2 );
not ( w1847 , w299 );
and ( w1848 , w1847 , g7 );
and ( w1849 , w1848 , g5 );
nor ( w1850 , w1588 , g1 );
nor ( w1851 , w1849 , w1850 );
and ( w1852 , w1851 , g4 );
nor ( w1853 , w1852 , g3 );
nor ( w1854 , w1853 , g3 );
nor ( w1855 , w1854 , w1395 );
and ( w1856 , w1855 , w8765 );
nor ( w1857 , w1856 , g9 );
nor ( w1858 , w1857 , g2 );
nor ( w1859 , w1858 , g2 );
and ( w1860 , w1859 , w8728 );
nor ( w1861 , w1846 , w1860 );
nor ( w1862 , w1861 , g9 );
and ( w1863 , w1862 , w8728 );
and ( w1864 , w1863 , w8735 );
nor ( w1865 , w1845 , w1864 );
and ( w1866 , w1865 , w8837 );
not ( w1867 , w1866 );
and ( w1868 , w1867 , w1608 );
and ( w1869 , w1802 , w8792 );
not ( w1870 , w1869 );
and ( w1871 , w1870 , w1567 );
and ( w1872 , w1871 , w8845 );
nor ( w1873 , w1868 , w1872 );
and ( w1874 , w1873 , w7934 );
nor ( w1875 , w1874 , g1 );
nor ( w1876 , w1875 , g1 );
not ( w1877 , w1876 );
and ( w1878 , w1877 , w1567 );
and ( w1879 , w1878 , w8735 );
and ( w1880 , w1879 , w8728 );
nor ( w1881 , w1880 , w1778 );
nor ( w1882 , w1881 , g7 );
and ( w1883 , w1882 , w8845 );
nor ( w1884 , w1883 , g13 );
not ( w1885 , w1884 );
and ( w1886 , w1885 , w1751 );
nor ( w1887 , w1886 , g16 );
not ( w1888 , w1843 );
and ( w1889 , w1888 , w1887 );
nor ( w1890 , w1889 , g6 );
and ( w1891 , w1890 , w8735 );
nor ( w1892 , w1891 , g13 );
not ( w1893 , w1892 );
and ( w1894 , w1893 , w1751 );
nor ( w1895 , w1894 , g16 );
not ( w1896 , w1640 );
and ( w1897 , w1896 , w1895 );
and ( w1898 , w92 , g4 );
and ( w1899 , w1898 , g2 );
nor ( w1900 , w1899 , g10 );
and ( w1901 , w1900 , g4 );
nor ( w1902 , w1897 , w1901 );
and ( w1903 , w1902 , g12 );
nor ( w1904 , w1903 , w1829 );
and ( w1905 , w1904 , w1950 );
nor ( w1906 , w1905 , g3 );
and ( w1907 , w1906 , w408 );
and ( w1908 , w1907 , g2 );
nor ( w1909 , w1908 , w1795 );
and ( w1910 , w1909 , w1838 );
not ( w1911 , w1910 );
and ( w1912 , w1911 , w1567 );
nor ( w1913 , w1912 , g1 );
nor ( w1914 , w1913 , g3 );
and ( w1915 , w1914 , g7 );
not ( w1916 , w1915 );
and ( w1917 , w1916 , w1887 );
nor ( w1918 , w1917 , g6 );
and ( w1919 , w1918 , w8735 );
nor ( w1920 , w1919 , g13 );
not ( w1921 , w1920 );
and ( w1922 , w1921 , w1751 );
nor ( w1923 , w1922 , g16 );
not ( w1924 , w1633 );
and ( w1925 , w1924 , w1923 );
and ( w1926 , w1925 , w1948 );
and ( w1927 , w1926 , w1950 );
nor ( w1928 , w1927 , g9 );
and ( w1929 , w1928 , g2 );
nor ( w1930 , w1929 , w1795 );
and ( w1931 , w1930 , w1838 );
not ( w1932 , w1931 );
and ( w1933 , w1932 , w1567 );
and ( w1934 , w1933 , w8792 );
nor ( w1935 , w1934 , g1 );
nor ( w1936 , w1935 , g3 );
and ( w1937 , w1936 , g7 );
not ( w1938 , w1937 );
and ( w1939 , w1938 , w1887 );
nor ( w1940 , w1939 , g6 );
and ( w1941 , w1940 , w8735 );
nor ( w1942 , w1941 , g13 );
not ( w1943 , w1942 );
and ( w1944 , w1943 , w1751 );
nor ( w1945 , w1944 , g16 );
not ( w1946 , w1604 );
and ( w1947 , w1946 , w1945 );
not ( w1948 , w1829 );
and ( w1949 , w1947 , w1948 );
not ( w1950 , w1824 );
and ( w1951 , w1949 , w1950 );
nor ( w1952 , w1951 , g9 );
and ( w1953 , w1952 , g2 );
nor ( w1954 , w1953 , w1795 );
and ( w1955 , w1954 , w1838 );
not ( w1956 , w1955 );
and ( w1957 , w1956 , w1567 );
and ( w1958 , w1957 , w8792 );
nor ( w1959 , w1958 , g1 );
nor ( w1960 , w1959 , g3 );
and ( w1961 , w1960 , g7 );
not ( w1962 , w1961 );
and ( w1963 , w1962 , w1887 );
nor ( w1964 , w1963 , g6 );
and ( w1965 , w1964 , w8735 );
nor ( w1966 , w1965 , g13 );
not ( w1967 , w1966 );
and ( w1968 , w1967 , w1751 );
nor ( w1969 , w1968 , g16 );
and ( w1970 , w6851 , w1969 );
and ( w1971 , g4 , g6 );
not ( w1972 , w1971 );
and ( w1973 , w1970 , w1972 );
nor ( w1974 , w1973 , g1 );
and ( w1975 , w1974 , g4 );
and ( w1976 , w1975 , w1751 );
not ( w1977 , w1976 );
and ( w1978 , w1588 , w1977 );
not ( w1979 , w1978 );
and ( w1980 , w1979 , g4 );
nor ( w1981 , w27 , g4 );
nor ( w1982 , w1981 , g9 );
nor ( w1983 , w1982 , g1 );
and ( w1984 , w8742 , g3 );
and ( w1985 , w1984 , w8769 );
nor ( w1986 , w1985 , g5 );
and ( w1987 , w1986 , w8742 );
nor ( w1988 , w1987 , g2 );
nor ( w1989 , w1988 , g2 );
nor ( w1990 , w1989 , g4 );
and ( w1991 , w1990 , w8765 );
nor ( w1992 , w1991 , g9 );
and ( w1993 , w8769 , w1244 );
nor ( w1994 , w1993 , g5 );
and ( w1995 , w1994 , w8742 );
not ( w1996 , w1995 );
and ( w1997 , w1996 , g2 );
not ( w1998 , w1997 );
and ( w1999 , w1998 , g2 );
nor ( w2000 , w1999 , g1 );
and ( w2001 , w2000 , w8765 );
and ( w2002 , w2001 , w8860 );
and ( w2003 , w2002 , w8765 );
and ( w2004 , w2003 , w8860 );
nor ( w2005 , w1430 , w2004 );
nor ( w2006 , w1992 , w2005 );
and ( w2007 , w2006 , g6 );
and ( w2008 , w2007 , w526 );
nor ( w2009 , w1982 , g9 );
nor ( w2010 , w2009 , g1 );
nor ( w2011 , w2010 , g1 );
nor ( w2012 , w2011 , g6 );
nor ( w2013 , w2012 , g6 );
nor ( w2014 , w2013 , g9 );
nor ( w2015 , w2014 , g6 );
and ( w2016 , w2015 , w8792 );
and ( w2017 , w2016 , g3 );
nor ( w2018 , w2008 , w2017 );
nor ( w2019 , w2018 , g4 );
nor ( w2020 , g1 , w663 );
and ( w2021 , w2020 , g2 );
and ( w2022 , w1516 , w7783 );
nor ( w2023 , w2021 , w2022 );
not ( w2024 , w2023 );
and ( w2025 , w2024 , g6 );
and ( w2026 , w2025 , w8860 );
and ( w2027 , w2026 , w361 );
nor ( w2028 , w2027 , g1 );
not ( w2029 , w2028 );
and ( w2030 , w2029 , g6 );
and ( w2031 , w2030 , w8735 );
and ( w2032 , w2031 , w8860 );
and ( w2033 , w2032 , w1751 );
nor ( w2034 , w1430 , w2033 );
and ( w2035 , w2034 , w8792 );
not ( w2036 , w770 );
and ( w2037 , w2036 , g6 );
not ( w2038 , w2037 );
and ( w2039 , w2038 , g6 );
not ( w2040 , w2035 );
and ( w2041 , w2040 , w2039 );
and ( w2042 , w2041 , w8860 );
not ( w2043 , w2042 );
and ( w2044 , w2043 , w1969 );
not ( w2045 , w2044 );
and ( w2046 , w2045 , w1567 );
and ( w2047 , w2046 , w8860 );
nor ( w2048 , w2019 , w2047 );
not ( w2049 , w2048 );
and ( w2050 , w2049 , w1751 );
and ( w2051 , w1983 , w2050 );
nor ( w2052 , w2051 , g1 );
not ( w2053 , w2052 );
and ( w2054 , w2053 , g3 );
nor ( w2055 , w2054 , w2047 );
nor ( w2056 , w2055 , g4 );
nor ( w2057 , w1980 , w2056 );
and ( w2058 , w1586 , w2148 );
nor ( w2059 , w2058 , g10 );
not ( w2060 , w2059 );
and ( w2061 , w2060 , g9 );
nor ( w2062 , w2061 , w471 );
nor ( w2063 , w2062 , g3 );
and ( w2064 , w2063 , g5 );
and ( w2065 , w512 , g7 );
and ( w2066 , w512 , w8742 );
and ( w2067 , w2066 , w59 );
nor ( w2068 , w2065 , w2067 );
not ( w2069 , w2068 );
and ( w2070 , w2069 , w17 );
and ( w2071 , w2070 , w2148 );
nor ( w2072 , g9 , w2071 );
and ( w2073 , w73 , w8769 );
not ( w2074 , w2073 );
and ( w2075 , w2074 , g10 );
nor ( w2076 , w2075 , g7 );
nor ( w2077 , w2076 , g7 );
not ( w2078 , w2077 );
and ( w2079 , w2078 , g8 );
not ( w2080 , w2079 );
and ( w2081 , w2080 , g8 );
nor ( w2082 , w2072 , w2081 );
not ( w2083 , w1582 );
and ( w2084 , w1521 , w2083 );
and ( w2085 , w2084 , g9 );
and ( w2086 , w2085 , w7783 );
nor ( w2087 , w2086 , w2071 );
nor ( w2088 , w2087 , g2 );
and ( w2089 , w2088 , w8845 );
and ( w2090 , w2089 , w8735 );
and ( w2091 , w2090 , w2148 );
and ( w2092 , w2082 , w2091 );
and ( w2093 , w2092 , w8769 );
nor ( w2094 , w2064 , w2093 );
nor ( w2095 , w566 , g5 );
and ( w2096 , w2095 , w8765 );
and ( w2097 , w2096 , g10 );
nor ( w2098 , w2097 , g7 );
nor ( w2099 , w2098 , g7 );
not ( w2100 , w2099 );
and ( w2101 , w2100 , g8 );
not ( w2102 , w2101 );
and ( w2103 , w2102 , g8 );
not ( w2104 , w2103 );
and ( w2105 , w2104 , w1844 );
and ( w2106 , w2105 , w27 );
and ( w2107 , w2106 , w8845 );
not ( w2108 , w2094 );
and ( w2109 , w2108 , w2107 );
and ( w2110 , w2109 , w8792 );
and ( w2111 , w2110 , w2148 );
nor ( w2112 , w1572 , w2111 );
not ( w2113 , w2112 );
and ( w2114 , w2113 , w27 );
and ( w2115 , w59 , g10 );
nor ( w2116 , w2115 , g7 );
nor ( w2117 , w2116 , g3 );
nor ( w2118 , w2117 , g5 );
nor ( w2119 , w2118 , g3 );
and ( w2120 , w2119 , w8860 );
and ( w2121 , w2120 , w8765 );
and ( w2122 , w2121 , w8845 );
and ( w2123 , w2122 , w8792 );
and ( w2124 , w2123 , g10 );
and ( w2125 , w2124 , g8 );
and ( w2126 , w2125 , w59 );
nor ( w2127 , w2126 , g5 );
and ( w2128 , w2127 , w8765 );
and ( w2129 , w2128 , w8735 );
and ( w2130 , w2129 , w8792 );
and ( w2131 , w2130 , g10 );
nor ( w2132 , w2131 , g7 );
and ( w2133 , w2132 , w8845 );
nor ( w2134 , w2133 , g7 );
not ( w2135 , w2134 );
and ( w2136 , w2135 , g8 );
not ( w2137 , w2136 );
and ( w2138 , w2137 , g8 );
nor ( w2139 , w2138 , g6 );
and ( w2140 , w2114 , w2139 );
and ( w2141 , w2140 , w2148 );
nor ( w2142 , w2141 , g3 );
and ( w2143 , w2142 , w8860 );
and ( w2144 , w2143 , w8792 );
not ( w2145 , w2144 );
and ( w2146 , w2145 , w1567 );
and ( w2147 , w2146 , w8845 );
not ( w2148 , w2057 );
and ( w2149 , w2147 , w2148 );
not ( w2150 , w1535 );
and ( w2151 , w2150 , w2149 );
and ( w2152 , w2151 , g3 );
not ( w2153 , w2152 );
and ( w2154 , w2153 , g13 );
not ( w2155 , w2154 );
and ( w2156 , w2155 , g3 );
and ( w2157 , w1521 , w400 );
and ( w2158 , w1531 , w8735 );
nor ( w2159 , w2157 , w2158 );
and ( w2160 , w2159 , g14 );
and ( w2161 , w2160 , w8168 );
nor ( w2162 , w2161 , g1 );
not ( w2163 , w2162 );
and ( w2164 , w2163 , g11 );
and ( w2165 , w1527 , g2 );
nor ( w2166 , w2165 , w2158 );
and ( w2167 , w2166 , w8837 );
nor ( w2168 , w2167 , g3 );
and ( w2169 , w2168 , w8792 );
not ( w2170 , w2164 );
and ( w2171 , w2170 , w2169 );
and ( w2172 , w2171 , w8845 );
not ( w2173 , w2172 );
and ( w2174 , w2173 , g16 );
not ( w2175 , w2174 );
and ( w2176 , w2175 , w2149 );
and ( w2177 , w77 , w27 );
and ( w2178 , w2177 , w33 );
nor ( w2179 , w2178 , g5 );
and ( w2180 , w2179 , w8765 );
and ( w2181 , w2180 , w8860 );
and ( w2182 , w2181 , g10 );
not ( w2183 , w2182 );
and ( w2184 , w2183 , g8 );
nor ( w2185 , w2184 , g7 );
and ( w2186 , w2185 , g8 );
not ( w2187 , w2186 );
and ( w2188 , w2176 , w2187 );
and ( w2189 , w77 , g8 );
nor ( w2190 , g4 , g9 );
and ( w2191 , w2189 , w2190 );
and ( w2192 , w2191 , g10 );
nor ( w2193 , w2192 , g5 );
and ( w2194 , w2193 , w8765 );
and ( w2195 , w2194 , w8860 );
and ( w2196 , w2195 , g10 );
nor ( w2197 , w2196 , g7 );
and ( w2198 , w2197 , w8735 );
nor ( w2199 , w2198 , g7 );
not ( w2200 , w2199 );
and ( w2201 , w2200 , g8 );
not ( w2202 , w2201 );
and ( w2203 , w2202 , g8 );
not ( w2204 , w2203 );
and ( w2205 , w2204 , w2149 );
and ( w2206 , w2205 , w8735 );
and ( w2207 , w2188 , w2206 );
nor ( w2208 , g2 , w2081 );
and ( w2209 , w2208 , w8742 );
and ( w2210 , w2209 , w8769 );
and ( w2211 , w2210 , g8 );
and ( w2212 , w2211 , w1844 );
and ( w2213 , w2212 , w2190 );
nor ( w2214 , w2213 , g5 );
and ( w2215 , w2214 , w8860 );
nor ( w2216 , w2215 , g3 );
nor ( w2217 , w2216 , g7 );
and ( w2218 , w2217 , g8 );
nor ( w2219 , w2218 , g2 );
nor ( w2220 , w2219 , g9 );
not ( w2221 , w400 );
and ( w2222 , w2221 , w2220 );
nor ( w2223 , w2222 , g1 );
nor ( w2224 , g9 , g6 );
and ( w2225 , w2224 , w1567 );
and ( w2226 , w2223 , w2225 );
and ( w2227 , w2226 , w361 );
nor ( w2228 , w2227 , g9 );
nor ( w2229 , w2228 , g3 );
and ( w2230 , w2229 , w8845 );
and ( w2231 , w2230 , w8792 );
and ( w2232 , w2207 , w2231 );
and ( w2233 , w2232 , g4 );
and ( w2234 , w2233 , w8742 );
and ( w2235 , w2107 , w8828 );
and ( w2236 , w2235 , g10 );
nor ( w2237 , w2236 , g11 );
and ( w2238 , w2237 , w8819 );
and ( w2239 , w2238 , g10 );
and ( w2240 , w2239 , w8168 );
not ( w2241 , w2240 );
and ( w2242 , w2241 , w2225 );
not ( w2243 , w2242 );
and ( w2244 , w2243 , g14 );
nor ( w2245 , w2244 , g5 );
and ( w2246 , w2245 , w7783 );
nor ( w2247 , w2246 , g9 );
and ( w2248 , w2247 , w8769 );
nor ( w2249 , w2248 , g7 );
nor ( w2250 , w2249 , g2 );
and ( w2251 , w2250 , w8742 );
nor ( w2252 , w2251 , g4 );
not ( w2253 , w2252 );
and ( w2254 , w2253 , g12 );
not ( w2255 , w2254 );
and ( w2256 , w2255 , g8 );
nor ( w2257 , w2256 , g4 );
and ( w2258 , w2257 , g8 );
nor ( w2259 , w2157 , w1531 );
not ( w2260 , w2259 );
and ( w2261 , w2260 , g9 );
nor ( w2262 , w1235 , g7 );
and ( w2263 , w2262 , w8769 );
and ( w2264 , w27 , w2263 );
nor ( w2265 , w2264 , g7 );
and ( w2266 , w2265 , w8860 );
and ( w2267 , w2266 , w8769 );
not ( w2268 , w2267 );
and ( w2269 , w2268 , g10 );
and ( w2270 , w2269 , w8767 );
nor ( w2271 , w2270 , g8 );
nor ( w2272 , w2271 , g1 );
and ( w2273 , w2272 , w1347 );
and ( w2274 , w2273 , w8765 );
and ( w2275 , w2274 , w8735 );
not ( w2276 , w2275 );
and ( w2277 , w2276 , g11 );
and ( w2278 , w2277 , g14 );
and ( w2279 , w2278 , w8168 );
and ( w2280 , w2279 , g13 );
nor ( w2281 , w2280 , g6 );
not ( w2282 , w2281 );
and ( w2283 , w2282 , g16 );
nor ( w2284 , w2283 , g3 );
and ( w2285 , w2284 , w8845 );
and ( w2286 , w2285 , w1567 );
and ( w2287 , w2286 , w8792 );
and ( w2288 , w2287 , g10 );
and ( w2289 , w2288 , g2 );
and ( w2290 , w42 , w1567 );
and ( w2291 , w2290 , g7 );
and ( w2292 , w2291 , g4 );
and ( w2293 , w44 , w2149 );
nor ( w2294 , w2292 , w2293 );
and ( w2295 , w408 , g4 );
and ( w2296 , w44 , w17 );
nor ( w2297 , w2296 , w1786 );
not ( w2298 , w2297 );
and ( w2299 , w2298 , g15 );
nor ( w2300 , w2299 , w1648 );
not ( w2301 , w2300 );
and ( w2302 , w2301 , w2149 );
and ( w2303 , w2302 , w8792 );
and ( w2304 , w2303 , w361 );
and ( w2305 , w2304 , w7783 );
nor ( w2306 , w2295 , w2305 );
not ( w2307 , w2306 );
and ( w2308 , w2307 , w2149 );
and ( w2309 , w2308 , w7783 );
and ( w2310 , w2309 , w2231 );
not ( w2311 , w2294 );
and ( w2312 , w2311 , w2310 );
nor ( w2313 , w2289 , w2312 );
nor ( w2314 , w2313 , g9 );
not ( w2315 , w2314 );
and ( w2316 , w2315 , g11 );
and ( w2317 , w2316 , g14 );
and ( w2318 , w2317 , w8168 );
and ( w2319 , w2318 , g13 );
nor ( w2320 , w2319 , g1 );
and ( w2321 , w2320 , w8845 );
not ( w2322 , w2321 );
and ( w2323 , w2322 , g16 );
and ( w2324 , w1569 , w27 );
nor ( w2325 , w2324 , g4 );
not ( w2326 , w2325 );
and ( w2327 , w2326 , g2 );
nor ( w2328 , g9 , w2310 );
nor ( w2329 , w2328 , g6 );
and ( w2330 , w2329 , w7783 );
and ( w2331 , w2330 , w2149 );
and ( w2332 , w2331 , w2206 );
and ( w2333 , w2332 , w2231 );
nor ( w2334 , w2327 , w2333 );
not ( w2335 , w2334 );
and ( w2336 , w2335 , w2149 );
and ( w2337 , w2336 , w8735 );
and ( w2338 , w2337 , w8792 );
and ( w2339 , w2338 , w361 );
and ( w2340 , w2339 , g2 );
nor ( w2341 , w2340 , w2333 );
and ( w2342 , w8765 , w2341 );
not ( w2343 , w2342 );
and ( w2344 , w2343 , g2 );
nor ( w2345 , w2344 , w2333 );
not ( w2346 , w2345 );
and ( w2347 , w2346 , w2149 );
and ( w2348 , w2347 , w8735 );
and ( w2349 , w2348 , w8792 );
not ( w2350 , w2323 );
and ( w2351 , w2350 , w2349 );
and ( w2352 , g4 , w8742 );
and ( w2353 , w2351 , w2401 );
nor ( w2354 , w2261 , w2353 );
nor ( w2355 , w2293 , g2 );
not ( w2356 , w2355 );
and ( w2357 , w2356 , g10 );
and ( w2358 , w2312 , w8730 );
not ( w2359 , w2358 );
and ( w2360 , w2359 , g12 );
and ( w2361 , w2360 , g16 );
not ( w2362 , w2361 );
and ( w2363 , w2362 , w2349 );
and ( w2364 , w2363 , w2401 );
nor ( w2365 , w2357 , w2364 );
and ( w2366 , w2365 , g12 );
and ( w2367 , w2366 , w8837 );
and ( w2368 , w2367 , g14 );
and ( w2369 , w2368 , w8168 );
and ( w2370 , w2369 , g13 );
nor ( w2371 , w2370 , g6 );
not ( w2372 , w2371 );
and ( w2373 , w2372 , g16 );
not ( w2374 , w2373 );
and ( w2375 , w2374 , w2349 );
and ( w2376 , w2375 , w2401 );
and ( w2377 , g12 , w2376 );
nor ( w2378 , w2377 , g10 );
not ( w2379 , w2378 );
and ( w2380 , w2379 , g2 );
nor ( w2381 , w2380 , w2312 );
and ( w2382 , g10 , g2 );
nor ( w2383 , w2382 , w1531 );
not ( w2384 , w2383 );
and ( w2385 , w2384 , g9 );
nor ( w2386 , w2385 , g11 );
and ( w2387 , w2386 , g14 );
and ( w2388 , w2387 , w8168 );
nor ( w2389 , w2388 , g1 );
not ( w2390 , w2389 );
and ( w2391 , w2381 , w2390 );
and ( w2392 , w2391 , w8837 );
and ( w2393 , w2392 , g14 );
and ( w2394 , w2393 , g13 );
nor ( w2395 , w2394 , g1 );
and ( w2396 , w2395 , w8845 );
not ( w2397 , w2396 );
and ( w2398 , w2397 , g16 );
not ( w2399 , w2398 );
and ( w2400 , w2399 , w2349 );
not ( w2401 , w2352 );
and ( w2402 , w2400 , w2401 );
not ( w2403 , w2354 );
and ( w2404 , w2403 , w2402 );
not ( w2405 , w2258 );
and ( w2406 , w2405 , w2404 );
nor ( w2407 , w2234 , w2406 );
not ( w2408 , w2156 );
and ( w2409 , w2408 , w2407 );
nor ( w2410 , w2409 , g6 );
and ( w2411 , w2410 , w8792 );
nor ( w2412 , w1517 , w2411 );
nor ( w2413 , w2412 , g3 );
and ( w2414 , w2413 , g2 );
and ( w2415 , w2414 , w8767 );
and ( w2416 , w2415 , g6 );
nor ( w2417 , w2416 , w2411 );
nor ( w2418 , w1515 , w2417 );
and ( w2419 , w2418 , w8860 );
and ( w2420 , w2419 , w27 );
nor ( w2421 , w2420 , g4 );
nor ( w2422 , w2421 , w2412 );
and ( w2423 , w2422 , w8767 );
nor ( w2424 , w2423 , w1350 );
nor ( w2425 , w1414 , w33 );
nor ( w2426 , w2425 , g3 );
and ( w2427 , w2426 , w8742 );
and ( w2428 , w2427 , w8860 );
and ( w2429 , w2428 , w8767 );
nor ( w2430 , w2429 , g7 );
not ( w2431 , w2430 );
and ( w2432 , w2431 , w17 );
nor ( w2433 , w2432 , g4 );
and ( w2434 , w2433 , w8767 );
and ( w2435 , w2434 , w8769 );
nor ( w2436 , w2424 , w2435 );
and ( w2437 , w2436 , w8765 );
and ( w2438 , w2437 , w8792 );
and ( w2439 , w2438 , g2 );
and ( w2440 , w2439 , w361 );
and ( w2441 , w2440 , g6 );
nor ( w2442 , w2441 , w2411 );
and ( w2443 , w2590 , w2442 );
and ( w2444 , w1517 , g9 );
nor ( w2445 , w2444 , w2411 );
and ( w2446 , w2443 , w2445 );
not ( w2447 , w2446 );
and ( w2448 , w2447 , g2 );
and ( w2449 , w1552 , w1361 );
nor ( w2450 , w2449 , g10 );
nor ( w2451 , g10 , g11 );
nor ( w2452 , w2450 , w2451 );
and ( w2453 , w2452 , w8735 );
nor ( w2454 , w2453 , w122 );
and ( w2455 , w2454 , g14 );
not ( w2456 , w2455 );
and ( w2457 , w2456 , g6 );
nor ( w2458 , w2457 , w2411 );
nor ( w2459 , w2458 , g1 );
and ( w2460 , w2459 , w8735 );
and ( w2461 , w2460 , g6 );
nor ( w2462 , w2461 , w2411 );
not ( w2463 , w2462 );
and ( w2464 , w2463 , w1521 );
nor ( w2465 , w2464 , g12 );
and ( w2466 , w2459 , w1521 );
and ( w2467 , w2466 , g9 );
and ( w2468 , w8730 , g11 );
and ( w2469 , w1588 , w8769 );
and ( w2470 , w2469 , w8742 );
nor ( w2471 , w2470 , g11 );
and ( w2472 , w2471 , g13 );
and ( w2473 , w2472 , g16 );
not ( w2474 , w2473 );
and ( w2475 , w2474 , g6 );
nor ( w2476 , w2475 , w2411 );
nor ( w2477 , w2476 , g1 );
not ( w2478 , w2468 );
and ( w2479 , w2478 , w2477 );
and ( w2480 , w2479 , w408 );
not ( w2481 , w2480 );
and ( w2482 , w2481 , g13 );
and ( w2483 , w2482 , g16 );
not ( w2484 , w2483 );
and ( w2485 , w2484 , g6 );
nor ( w2486 , w2485 , w2411 );
nor ( w2487 , w2486 , g1 );
nor ( w2488 , w2467 , w2487 );
nor ( w2489 , w2488 , g3 );
nor ( w2490 , w2489 , w122 );
and ( w2491 , w2490 , g13 );
and ( w2492 , w2491 , g14 );
and ( w2493 , w2492 , g16 );
not ( w2494 , w2493 );
and ( w2495 , w2494 , g6 );
nor ( w2496 , w2495 , w2411 );
nor ( w2497 , w2496 , g1 );
and ( w2498 , w2466 , g4 );
nor ( w2499 , w2498 , w27 );
and ( w2500 , w2499 , w8168 );
and ( w2501 , w2500 , g13 );
and ( w2502 , w2501 , g14 );
not ( w2503 , w2502 );
and ( w2504 , w2503 , g6 );
nor ( w2505 , w2504 , w2411 );
nor ( w2506 , w2505 , g1 );
and ( w2507 , w2497 , w2506 );
and ( w2508 , w8792 , g4 );
nor ( w2509 , w2508 , w27 );
not ( w2510 , w2509 );
and ( w2511 , w2510 , g6 );
nor ( w2512 , w2511 , w2411 );
nor ( w2513 , w2512 , g1 );
and ( w2514 , w2513 , w33 );
not ( w2515 , w2514 );
and ( w2516 , w2515 , g10 );
nor ( w2517 , w2516 , g3 );
and ( w2518 , w2517 , g6 );
nor ( w2519 , w2518 , w2411 );
nor ( w2520 , w2519 , g1 );
and ( w2521 , w2507 , w2520 );
and ( w2522 , w2521 , w8735 );
nor ( w2523 , w2522 , w122 );
and ( w2524 , w2523 , g13 );
and ( w2525 , w2524 , g14 );
and ( w2526 , w2525 , g16 );
not ( w2527 , w2526 );
and ( w2528 , w2527 , g6 );
nor ( w2529 , w2528 , w2411 );
nor ( w2530 , w2529 , g1 );
not ( w2531 , w2465 );
and ( w2532 , w2531 , w2530 );
nor ( w2533 , w2532 , w122 );
and ( w2534 , w2533 , g13 );
and ( w2535 , w2534 , g14 );
and ( w2536 , w2535 , g16 );
not ( w2537 , w2536 );
and ( w2538 , w2537 , g6 );
nor ( w2539 , w2538 , w2411 );
nor ( w2540 , w2539 , g1 );
and ( w2541 , w2540 , w8735 );
nor ( w2542 , w33 , w1361 );
nor ( w2543 , w2542 , g1 );
and ( w2544 , w8792 , g8 );
not ( w2545 , w2544 );
and ( w2546 , w2545 , g8 );
not ( w2547 , w2546 );
and ( w2548 , w2547 , g9 );
not ( w2549 , w2548 );
and ( w2550 , w2549 , w765 );
not ( w2551 , w2550 );
and ( w2552 , w2551 , g6 );
nor ( w2553 , w2552 , w2411 );
nor ( w2554 , w2553 , g1 );
and ( w2555 , w2543 , w2554 );
not ( w2556 , w2451 );
and ( w2557 , w2555 , w2556 );
nor ( w2558 , w2557 , w122 );
and ( w2559 , w2558 , g14 );
not ( w2560 , w2559 );
and ( w2561 , w2560 , g6 );
nor ( w2562 , w2561 , w2411 );
nor ( w2563 , w2562 , g1 );
and ( w2564 , w2563 , w1521 );
and ( w2565 , w2564 , g3 );
nor ( w2566 , w2565 , w122 );
and ( w2567 , w2566 , g13 );
and ( w2568 , w2567 , g14 );
not ( w2569 , w2568 );
and ( w2570 , w2569 , g6 );
nor ( w2571 , w2570 , w2411 );
nor ( w2572 , w2571 , g1 );
nor ( w2573 , w2541 , w2572 );
and ( w2574 , w2573 , w8168 );
and ( w2575 , w2574 , g13 );
and ( w2576 , w2575 , g14 );
and ( w2577 , w2576 , g16 );
not ( w2578 , w2577 );
and ( w2579 , w2578 , g6 );
nor ( w2580 , w2579 , w2411 );
nor ( w2581 , w2580 , g1 );
not ( w2582 , w2581 );
and ( w2583 , w2582 , g13 );
and ( w2584 , w2583 , g16 );
and ( w2585 , g6 , g2 );
and ( w2586 , w2413 , w2585 );
nor ( w2587 , w2022 , w2411 );
not ( w2588 , w2586 );
and ( w2589 , w2588 , w2587 );
not ( w2590 , w1514 );
and ( w2591 , w2590 , w2589 );
not ( w2592 , w2591 );
and ( w2593 , w2592 , w1751 );
and ( w2594 , w2593 , g6 );
nor ( w2595 , w2594 , w2411 );
nor ( w2596 , w2584 , w2595 );
and ( w2597 , w2022 , w2596 );
nor ( w2598 , w2597 , w2411 );
not ( w2599 , w2448 );
and ( w2600 , w2599 , w2598 );
nor ( w2601 , w2600 , w2595 );
nor ( w2602 , w2601 , g1 );
not ( w2603 , w2602 );
and ( w2604 , w2603 , g10 );
not ( w2605 , w2604 );
and ( w2606 , w2605 , g10 );
nor ( w2607 , g7 , g12 );
nor ( w2608 , w1421 , g9 );
and ( w2609 , w2608 , w8860 );
nor ( w2610 , w2609 , g3 );
not ( w2611 , w2607 );
and ( w2612 , w2611 , w2610 );
nor ( w2613 , w2612 , g1 );
nor ( w2614 , w2613 , g3 );
nor ( w2615 , w2614 , g2 );
and ( w2616 , w2615 , w8730 );
nor ( w2617 , w2616 , g10 );
and ( w2618 , w2617 , w7783 );
and ( w2619 , g6 , w8765 );
not ( w2620 , w2618 );
and ( w2621 , w2620 , w2619 );
and ( w2622 , w2621 , w408 );
nor ( w2623 , w2622 , g9 );
nor ( w2624 , w2623 , w2602 );
nor ( w2625 , w2624 , g16 );
nor ( w2626 , w2625 , w2602 );
nor ( w2627 , w2626 , w381 );
and ( w2628 , w2627 , g11 );
not ( w2629 , w2628 );
and ( w2630 , w2629 , g6 );
not ( w2631 , w1668 );
and ( w2632 , w2631 , w1567 );
nor ( w2633 , w2632 , g16 );
and ( w2634 , w2633 , g13 );
not ( w2635 , w2634 );
and ( w2636 , w2635 , w1567 );
nor ( w2637 , w2636 , w122 );
not ( w2638 , w2637 );
and ( w2639 , w2638 , w2601 );
nor ( w2640 , w2639 , g16 );
and ( w2641 , w2640 , g11 );
not ( w2642 , w2641 );
and ( w2643 , w2642 , w2601 );
and ( w2644 , w2643 , g6 );
nor ( w2645 , w2644 , w2411 );
not ( w2646 , w2645 );
and ( w2647 , w2630 , w2646 );
nor ( w2648 , w2647 , g1 );
and ( w2649 , w2648 , g13 );
nor ( w2650 , w2602 , w2649 );
nor ( w2651 , w2650 , g14 );
and ( w2652 , w2651 , w8168 );
nor ( w2653 , w2652 , w2602 );
not ( w2654 , w2653 );
and ( w2655 , w2654 , g11 );
not ( w2656 , w2655 );
and ( w2657 , w2656 , g6 );
nor ( w2658 , w2657 , g1 );
and ( w2659 , w2658 , g13 );
nor ( w2660 , w2606 , w2659 );
and ( w2661 , w2645 , w8792 );
not ( w2662 , w2661 );
and ( w2663 , w2660 , w2662 );
and ( w2664 , w2663 , g6 );
nor ( w2665 , w2411 , g1 );
not ( w2666 , w2664 );
and ( t_4 , w2666 , w2665 );
and ( w2667 , g2 , w8837 );
nor ( w2668 , g11 , w2667 );
nor ( w2669 , w2668 , g6 );
and ( w2670 , w7186 , g2 );
and ( w2671 , w2670 , g13 );
and ( w2672 , w2671 , w8828 );
and ( w2673 , w2672 , w8837 );
and ( w2674 , w2673 , w8765 );
and ( w2675 , w2674 , g1 );
nor ( w2676 , w381 , w1244 );
nor ( w2677 , w2676 , g9 );
nor ( w2678 , w2677 , w381 );
nor ( w2679 , w2678 , g1 );
and ( w2680 , w2679 , w8769 );
nor ( w2681 , w2680 , g5 );
nor ( w2682 , w2681 , w1987 );
and ( w2683 , w2682 , g6 );
and ( w2684 , w2683 , g3 );
and ( w2685 , w2684 , w8765 );
and ( w2686 , w2685 , w8860 );
nor ( w2687 , g4 , g1 );
and ( w2688 , w2686 , w2687 );
not ( w2689 , w2688 );
and ( w2690 , w2689 , g6 );
not ( w2691 , w2690 );
and ( w2692 , w2691 , g3 );
and ( w2693 , w2692 , w8765 );
nor ( w2694 , w2693 , g12 );
not ( w2695 , w2694 );
and ( w2696 , w2695 , g2 );
not ( w2697 , w2696 );
and ( w2698 , w2697 , g11 );
and ( w2699 , w2698 , w8819 );
not ( w2700 , w2699 );
and ( w2701 , w2700 , g2 );
not ( w2702 , w2701 );
and ( w2703 , w2702 , g2 );
and ( w2704 , w2703 , w8792 );
nor ( w2705 , w2704 , g9 );
nor ( w2706 , w2705 , g9 );
and ( w2707 , w2706 , w8828 );
and ( w2708 , w8860 , w2707 );
not ( w2709 , w2708 );
and ( w2710 , w2709 , g3 );
and ( w2711 , w8742 , g2 );
and ( w2712 , w2711 , w8860 );
and ( w2713 , w2712 , g6 );
and ( w2714 , w2713 , g15 );
not ( w2715 , w2714 );
and ( w2716 , w2715 , g6 );
and ( w2717 , w2716 , w8742 );
and ( w2718 , w2717 , w8860 );
and ( w2719 , w2718 , w8168 );
not ( w2720 , w2719 );
and ( w2721 , w2720 , w361 );
and ( w2722 , w2721 , g2 );
nor ( w2723 , w2710 , w2722 );
nor ( w2724 , g4 , g14 );
and ( w2725 , w2724 , w8168 );
and ( w2726 , w2725 , w8730 );
and ( w2727 , w2726 , g11 );
and ( w2728 , w8833 , g5 );
and ( w2729 , w2728 , w8728 );
and ( w2730 , w2729 , w8730 );
and ( w2731 , w2730 , g6 );
and ( w2732 , w2731 , g13 );
and ( w2733 , w2732 , g3 );
and ( w2734 , w2733 , w8828 );
and ( w2735 , w2734 , w8792 );
and ( w2736 , w2735 , w7141 );
and ( w2737 , w2736 , w8742 );
and ( w2738 , w2737 , g11 );
and ( w2739 , w2738 , w7783 );
nor ( w2740 , w2675 , w2739 );
not ( w2741 , w2740 );
and ( w2742 , w2741 , g14 );
nor ( w2743 , w2742 , w2739 );
not ( w2744 , w2727 );
and ( w2745 , w2744 , w2743 );
nor ( w2746 , g4 , g11 );
not ( w2747 , w2746 );
and ( w2748 , w2745 , w2747 );
nor ( w2749 , w2748 , g12 );
nor ( w2750 , w224 , w381 );
and ( w2751 , w2750 , g3 );
and ( w2752 , w2751 , g7 );
not ( w2753 , w2750 );
and ( w2754 , w2753 , g3 );
nor ( w2755 , w2754 , w1786 );
nor ( w2756 , w2754 , w381 );
and ( w2757 , w2756 , g11 );
and ( w2758 , w2757 , g13 );
and ( w2759 , w2758 , w7783 );
and ( w2760 , w2759 , w8792 );
and ( w2761 , w2760 , w8765 );
and ( w2762 , w2755 , w2761 );
and ( w2763 , w8742 , w2762 );
nor ( w2764 , w2752 , w2763 );
nor ( w2765 , g5 , g3 );
nor ( w2766 , w2764 , w2765 );
and ( w2767 , w2766 , g4 );
nor ( w2768 , w381 , g5 );
not ( w2769 , w2768 );
and ( w2770 , w2769 , g7 );
nor ( w2771 , w2770 , w381 );
and ( w2772 , w2771 , w8728 );
and ( w2773 , w7934 , g7 );
and ( w2774 , w2773 , g12 );
nor ( w2775 , w2772 , w2774 );
nor ( w2776 , w2775 , w59 );
not ( w2777 , w224 );
and ( w2778 , w2776 , w2777 );
and ( w2779 , w1707 , w7934 );
nor ( w2780 , w2778 , w2779 );
not ( w2781 , w2780 );
and ( w2782 , w2781 , g3 );
and ( w2783 , w7934 , g12 );
and ( w2784 , w2783 , w8735 );
nor ( w2785 , w2782 , w2784 );
nor ( w2786 , w2785 , g4 );
and ( w2787 , w2786 , g11 );
and ( w2788 , w2787 , g13 );
and ( w2789 , w2788 , w8792 );
and ( w2790 , w2789 , w8765 );
and ( w2791 , w2790 , w8828 );
nor ( w2792 , w2767 , w2791 );
not ( w2793 , w2792 );
and ( w2794 , w2793 , g11 );
and ( w2795 , w2794 , g6 );
and ( w2796 , w2795 , g13 );
and ( w2797 , w2784 , g4 );
and ( w2798 , w2797 , g11 );
and ( w2799 , w2798 , g6 );
and ( w2800 , w2799 , g13 );
and ( w2801 , w2800 , w7783 );
and ( w2802 , w2801 , w8792 );
and ( w2803 , w2802 , w8765 );
and ( w2804 , w2803 , w8828 );
nor ( w2805 , w2796 , w2804 );
nor ( w2806 , w2805 , g2 );
and ( w2807 , w2806 , w8792 );
and ( w2808 , w2807 , w8765 );
and ( w2809 , w2808 , w8828 );
not ( w2810 , w2809 );
and ( w2811 , w2743 , w2810 );
not ( w2812 , w2749 );
and ( w2813 , w2812 , w2811 );
and ( w2814 , w2813 , g6 );
and ( w2815 , w2814 , w8735 );
nor ( w2816 , w1852 , g12 );
and ( w2817 , w2816 , w8837 );
and ( w2818 , w2817 , g6 );
and ( w2819 , w2818 , w8735 );
nor ( w2820 , w2819 , g2 );
not ( w2821 , w2815 );
and ( w2822 , w2821 , w2820 );
and ( w2823 , w8728 , w59 );
and ( w2824 , w2823 , w8860 );
not ( w2825 , w2824 );
and ( w2826 , w2825 , g6 );
not ( w2827 , w2826 );
and ( w2828 , w2827 , w2743 );
and ( w2829 , w2824 , g6 );
and ( w2830 , g11 , w8845 );
nor ( w2831 , w2829 , w2830 );
not ( w2832 , w2831 );
and ( w2833 , w2832 , g3 );
nor ( w2834 , w2833 , g13 );
nor ( w2835 , w2834 , w2809 );
nor ( w2836 , w2835 , w381 );
and ( w2837 , w2836 , w7783 );
and ( w2838 , w2837 , w8792 );
and ( w2839 , w2838 , w8765 );
and ( w2840 , w2839 , w8828 );
not ( w2841 , w2840 );
and ( w2842 , w2828 , w2841 );
and ( w2843 , w2842 , g3 );
and ( w2844 , g6 , w8730 );
nor ( w2845 , w2844 , g10 );
not ( w2846 , w2845 );
and ( w2847 , w2846 , g6 );
nor ( w2848 , w2847 , g4 );
and ( w2849 , w2848 , w8837 );
and ( w2850 , w2849 , w8728 );
and ( w2851 , w2850 , w8735 );
nor ( w2852 , w2851 , g13 );
nor ( w2853 , w2852 , w2809 );
nor ( w2854 , w2853 , w381 );
and ( w2855 , w2854 , w7783 );
and ( w2856 , w2855 , w8792 );
and ( w2857 , w2856 , w8765 );
and ( w2858 , w2857 , w8828 );
not ( w2859 , w2843 );
and ( w2860 , w2859 , w2858 );
and ( w2861 , w2820 , w8819 );
nor ( w2862 , w2861 , w2809 );
nor ( w2863 , w2862 , w381 );
and ( w2864 , w2863 , w8792 );
and ( w2865 , w2864 , w8765 );
and ( w2866 , w2865 , w8828 );
and ( w2867 , w2860 , w2866 );
and ( w2868 , w2822 , w2867 );
not ( w2869 , w1244 );
and ( w2870 , w2869 , w2868 );
and ( w2871 , w2870 , g6 );
nor ( w2872 , w2871 , g3 );
not ( w2873 , w2872 );
and ( w2874 , w2873 , g11 );
nor ( w2875 , w2874 , w2809 );
not ( w2876 , w2875 );
and ( w2877 , w2876 , w2858 );
nor ( w2878 , w2877 , g3 );
nor ( w2879 , w2878 , g3 );
not ( w2880 , w2879 );
and ( w2881 , w2880 , w2811 );
and ( w2882 , w2881 , w7783 );
nor ( w2883 , w2882 , g2 );
nor ( w2884 , w2883 , g9 );
nor ( w2885 , w2884 , g9 );
nor ( w2886 , w2723 , w2885 );
and ( w2887 , w2886 , w289 );
not ( w2888 , w2887 );
and ( w2889 , w2888 , g2 );
nor ( w2890 , w2889 , w2885 );
nor ( w2891 , w2890 , g1 );
nor ( w2892 , w2891 , g9 );
nor ( w2893 , w2892 , g9 );
nor ( w2894 , w2675 , w2893 );
and ( w2895 , w2894 , w2743 );
nor ( w2896 , w1653 , w1613 );
and ( w2897 , w8223 , g17 );
and ( w2898 , w2897 , w8382 );
and ( w2899 , w2898 , g14 );
and ( w2900 , w2899 , w8860 );
and ( w2901 , w2900 , g10 );
and ( w2902 , w2901 , w7186 );
and ( w2903 , w2902 , g1 );
not ( w2904 , w2903 );
and ( w2905 , w2904 , w2894 );
not ( w2906 , w2905 );
and ( w2907 , w2906 , g13 );
and ( w2908 , w2907 , w8837 );
and ( w2909 , w2908 , g2 );
and ( w2910 , w2909 , g9 );
not ( w2911 , w2910 );
and ( w2912 , w2911 , w2894 );
nor ( w2913 , w2912 , g16 );
and ( w2914 , w2895 , g3 );
and ( w2915 , w2939 , g1 );
and ( w2916 , w2022 , g10 );
not ( w2917 , w2916 );
and ( w2918 , w2917 , g10 );
not ( w2919 , w2918 );
and ( w2920 , w2919 , w2895 );
and ( w2921 , w2920 , g8 );
not ( w2922 , w2921 );
and ( w2923 , w2922 , g8 );
not ( w2924 , w2923 );
and ( w2925 , w2924 , w2894 );
and ( w2926 , w2925 , w7783 );
nor ( w2927 , w2926 , g2 );
not ( w2928 , w2927 );
and ( w2929 , w2928 , g6 );
and ( w2930 , w2929 , w8792 );
and ( w2931 , w2930 , g9 );
not ( w2932 , w2931 );
and ( w2933 , w2932 , g9 );
not ( w2934 , w2933 );
and ( w2935 , w2934 , w2894 );
and ( w2936 , w2935 , w2895 );
not ( w2937 , w2739 );
and ( w2938 , w2937 , w381 );
not ( w2939 , w2742 );
and ( w2940 , w2938 , w2939 );
nor ( w2941 , w2940 , g2 );
and ( w2942 , w2941 , w8837 );
and ( w2943 , w2942 , g9 );
not ( w2944 , w2943 );
and ( w2945 , w2944 , w2894 );
nor ( w2946 , w2945 , g16 );
not ( w2947 , w2946 );
and ( w2948 , w2936 , w2947 );
and ( w2949 , w2948 , g6 );
not ( w2950 , w2949 );
and ( w2951 , w2950 , w2847 );
nor ( w2952 , w2951 , g1 );
not ( w2953 , w2952 );
and ( w2954 , w2953 , g13 );
and ( w2955 , w2954 , g12 );
not ( w2956 , w2955 );
and ( w2957 , w2956 , g9 );
not ( w2958 , w2957 );
and ( w2959 , w2958 , g9 );
not ( w2960 , w2959 );
and ( w2961 , w2960 , w2894 );
nor ( w2962 , w2961 , g16 );
not ( w2963 , w2915 );
and ( w2964 , w2963 , w2962 );
and ( w2965 , w2964 , g13 );
not ( w2966 , w2965 );
and ( w2967 , w2966 , w2894 );
and ( w2968 , w2967 , w2895 );
and ( w2969 , w2968 , w8735 );
not ( w2970 , w2969 );
and ( w2971 , w2970 , g12 );
not ( w2972 , w2971 );
and ( w2973 , w2972 , g9 );
not ( w2974 , w2973 );
and ( w2975 , w2974 , g9 );
not ( w2976 , w2975 );
and ( w2977 , w2976 , w2894 );
nor ( w2978 , w2977 , g16 );
not ( w2979 , w2914 );
and ( w2980 , w2979 , w2978 );
nor ( w2981 , w2913 , w2980 );
and ( w2982 , w2981 , w2895 );
and ( w2983 , w2982 , g3 );
not ( w2984 , w2983 );
and ( w2985 , w2984 , w2978 );
not ( w2986 , w2985 );
and ( w2987 , w2895 , w2986 );
and ( w2988 , w8828 , w2987 );
nor ( w2989 , w2988 , g5 );
and ( w2990 , w2989 , g7 );
nor ( w2991 , w2988 , g7 );
and ( w2992 , w2991 , w7070 );
nor ( w2993 , w2990 , w2992 );
not ( w2994 , w2993 );
and ( w2995 , w2994 , g17 );
and ( w2996 , w2995 , g12 );
and ( w2997 , w2996 , w8382 );
and ( w2998 , w2997 , g14 );
and ( w2999 , w2998 , g3 );
and ( w3000 , w2999 , g9 );
and ( w3001 , w3000 , w8860 );
and ( w3002 , w3001 , g13 );
and ( w3003 , w3002 , w8845 );
and ( w3004 , w3003 , w8730 );
not ( w3005 , w3004 );
and ( w3006 , w3005 , w2987 );
not ( w3007 , w3006 );
and ( w3008 , w3007 , g1 );
not ( w3009 , w3008 );
and ( w3010 , w3009 , w2987 );
not ( w3011 , w3010 );
and ( w3012 , w3011 , g2 );
not ( w3013 , w3012 );
and ( w3014 , w3013 , w2987 );
nor ( w3015 , w3014 , g11 );
not ( w3016 , w3015 );
nand ( t_5 , w3016 , w2987 );
nor ( w3017 , w2190 , g4 );
nor ( w3018 , w3017 , w79 );
nor ( w3019 , w3018 , g9 );
nor ( w3020 , w3019 , g5 );
and ( w3021 , w3020 , w8728 );
and ( w3022 , w3021 , g6 );
nor ( w3023 , g4 , w2687 );
nor ( w3024 , w3023 , g9 );
and ( w3025 , w3024 , g3 );
and ( w3026 , w3025 , w8769 );
nor ( w3027 , w3026 , g5 );
and ( w3028 , w1609 , w8728 );
and ( w3029 , w3028 , g6 );
nor ( w3030 , w3029 , g16 );
and ( w3031 , w3030 , g3 );
nor ( w3032 , g3 , g14 );
and ( w3033 , w3032 , w8730 );
and ( w3034 , w3033 , w8735 );
and ( w3035 , w3034 , g4 );
and ( w3036 , w3035 , w8742 );
and ( w3037 , g6 , w8828 );
and ( w3038 , w3037 , w8819 );
and ( w3039 , w3038 , g2 );
and ( w3040 , w3039 , w8792 );
and ( w3041 , w3040 , g7 );
nor ( w3042 , w3036 , w3041 );
and ( w3043 , w92 , w122 );
not ( w3044 , w3043 );
and ( w3045 , w3042 , w3044 );
and ( w3046 , w3045 , w7141 );
and ( w3047 , w3046 , w8730 );
not ( w3048 , w3047 );
and ( w3049 , w3048 , w3040 );
and ( w3050 , w3049 , w8728 );
and ( w3051 , w3050 , w8735 );
and ( w3052 , w3051 , g11 );
and ( w3053 , w3052 , w7997 );
and ( w3054 , w3040 , g12 );
and ( w3055 , w3054 , w8735 );
and ( w3056 , w3055 , g11 );
nor ( w3057 , w3053 , w3056 );
and ( w3058 , w244 , w8728 );
and ( w3059 , w3058 , w8828 );
and ( w3060 , w3059 , w8837 );
and ( w3061 , w3060 , w8819 );
nor ( w3062 , w467 , w3061 );
nor ( w3063 , w3062 , g12 );
and ( w3064 , w8845 , g12 );
and ( w3065 , w3064 , g2 );
nor ( w3066 , w3063 , w3065 );
nor ( w3067 , w3066 , g3 );
and ( w3068 , w3067 , w8828 );
and ( w3069 , w3068 , w8837 );
and ( w3070 , w3069 , w8819 );
and ( w3071 , w3070 , g2 );
and ( w3072 , w3071 , w8792 );
nor ( w3073 , w551 , g3 );
and ( w3074 , w3073 , w8819 );
and ( w3075 , w3074 , w8828 );
and ( w3076 , w3075 , w8765 );
nor ( w3077 , g11 , w3076 );
nor ( w3078 , w3077 , g3 );
and ( w3079 , w3078 , w8845 );
and ( w3080 , w3079 , w8819 );
and ( w3081 , w3080 , w8828 );
and ( w3082 , w3081 , w7997 );
and ( w3083 , w3082 , w7783 );
and ( w3084 , w3083 , w8765 );
nor ( w3085 , w3072 , w3084 );
nor ( w3086 , w3085 , w213 );
not ( w3087 , w3086 );
and ( w3088 , w3057 , w3087 );
nor ( w3089 , w3088 , w213 );
nor ( w3090 , w3031 , w3089 );
not ( w3091 , w3090 );
and ( w3092 , w3091 , g11 );
nor ( w3093 , w3092 , w3086 );
nor ( w3094 , w3093 , g13 );
and ( w3095 , w3094 , g2 );
nor ( w3096 , w3095 , w3084 );
nor ( w3097 , w3096 , w213 );
and ( w3098 , w3097 , w8792 );
not ( w3099 , w3027 );
and ( w3100 , w3099 , w3098 );
and ( w3101 , w3100 , g6 );
not ( w3102 , w3101 );
and ( w3103 , w3102 , g6 );
nor ( w3104 , w3103 , g16 );
and ( w3105 , w3104 , g3 );
nor ( w3106 , w3105 , w3089 );
not ( w3107 , w3106 );
and ( w3108 , w3107 , g11 );
nor ( w3109 , w3108 , w3086 );
nor ( w3110 , w3109 , g13 );
and ( w3111 , w3110 , g2 );
nor ( w3112 , w3111 , w3084 );
nor ( w3113 , w3112 , w213 );
and ( w3114 , w3113 , w8792 );
nor ( w3115 , w3114 , w3089 );
and ( w3116 , w3022 , w3115 );
not ( w3117 , w3116 );
and ( w3118 , w3117 , g3 );
nor ( w3119 , g6 , g12 );
nor ( w3120 , g14 , w122 );
and ( w3121 , w3120 , w8730 );
and ( w3122 , w299 , w3121 );
and ( w3123 , w3065 , w3491 );
and ( w3124 , w3123 , w8792 );
nor ( w3125 , w3119 , w3124 );
and ( w3126 , w8845 , w122 );
and ( w3127 , w3034 , g5 );
and ( w3128 , w3034 , w8742 );
nor ( w3129 , w3127 , w3128 );
and ( w3130 , w3129 , w3121 );
and ( w3131 , w5221 , g10 );
nor ( w3132 , w3130 , w3131 );
and ( w3133 , w3132 , g15 );
and ( w3134 , w3133 , w8845 );
and ( w3135 , w3134 , w8735 );
and ( w3136 , w3135 , w8819 );
and ( w3137 , w3136 , w7997 );
nor ( w3138 , w3126 , w3137 );
and ( w3139 , w3138 , w8728 );
nor ( w3140 , w3139 , g4 );
and ( w3141 , w3140 , w8735 );
and ( w3142 , w3141 , w8819 );
and ( w3143 , w3142 , w8828 );
and ( w3144 , w3143 , w7997 );
and ( w3145 , w3144 , w8792 );
nor ( w3146 , w3145 , g12 );
and ( w3147 , w3146 , w3115 );
nor ( w3148 , w3147 , g4 );
and ( w3149 , w3148 , w8735 );
and ( w3150 , w3149 , g11 );
nor ( w3151 , w3150 , w3086 );
nor ( w3152 , w3151 , g13 );
and ( w3153 , w3152 , w8828 );
and ( w3154 , w3153 , g2 );
and ( w3155 , w3154 , w7997 );
and ( w3156 , w3155 , w8792 );
nor ( w3157 , w3156 , w3084 );
and ( w3158 , w3115 , w3157 );
and ( w3159 , w3125 , w3158 );
not ( w3160 , w3159 );
and ( w3161 , w3160 , g4 );
not ( w3162 , w3161 );
and ( w3163 , w3162 , w3157 );
nor ( w3164 , w3163 , g3 );
and ( w3165 , w3164 , g11 );
nor ( w3166 , w3165 , w3086 );
nor ( w3167 , w3166 , g13 );
and ( w3168 , w3167 , w8828 );
and ( w3169 , w3168 , g2 );
and ( w3170 , w3169 , w7997 );
and ( w3171 , w3170 , w8792 );
nor ( w3172 , w3171 , w3084 );
not ( w3173 , w3118 );
and ( w3174 , w3173 , w3172 );
not ( w3175 , w3174 );
and ( w3176 , w3175 , g11 );
nor ( w3177 , w3176 , w3086 );
nor ( w3178 , w3177 , g13 );
and ( w3179 , w3178 , w8828 );
and ( w3180 , w3179 , g2 );
and ( w3181 , w3180 , w7997 );
and ( w3182 , w3181 , w8792 );
nor ( w3183 , w3182 , w3084 );
and ( w3184 , w473 , w8769 );
and ( w3185 , w3184 , w13 );
not ( w3186 , w3185 );
and ( w3187 , w3186 , g8 );
and ( w3188 , g10 , w6151 );
nor ( w3189 , w3188 , g7 );
and ( w3190 , w3189 , g10 );
not ( w3191 , w3190 );
and ( w3192 , w3191 , g10 );
nor ( w3193 , w3187 , w3192 );
and ( w3194 , w3193 , w17 );
and ( w3195 , w3194 , w27 );
and ( w3196 , w3195 , w8845 );
and ( w3197 , w3196 , w8792 );
and ( w3198 , w3197 , g10 );
nor ( w3199 , w3198 , w1786 );
nor ( w3200 , g3 , g6 );
not ( w3201 , w3199 );
and ( w3202 , w3201 , w3200 );
nor ( w3203 , w3202 , w270 );
and ( w3204 , w8728 , w3200 );
and ( w3205 , w770 , w5461 );
and ( w3206 , w3205 , w8730 );
and ( w3207 , w3206 , w17 );
nor ( w3208 , w3207 , w1786 );
not ( w3209 , w3208 );
and ( w3210 , w3209 , g12 );
and ( w3211 , w3210 , w8765 );
and ( w3212 , w3211 , g15 );
and ( w3213 , w3212 , g14 );
and ( w3214 , w27 , w3213 );
nor ( w3215 , w3204 , w3214 );
nor ( w3216 , w3215 , g7 );
nor ( w3217 , w3216 , w270 );
and ( w3218 , w3217 , w8860 );
nor ( w3219 , w3218 , g9 );
and ( w3220 , w3219 , w8845 );
and ( w3221 , w3220 , g15 );
and ( w3222 , w3221 , g14 );
and ( w3223 , w8735 , w3222 );
not ( w3224 , w3223 );
and ( w3225 , w3203 , w3224 );
and ( w3226 , w3225 , w8860 );
not ( w3227 , w3226 );
and ( w3228 , w3227 , g14 );
and ( w3229 , w3228 , g15 );
and ( w3230 , w3229 , w8845 );
and ( w3231 , w3230 , w8765 );
and ( w3232 , w8845 , g7 );
nor ( w3233 , w3232 , w1244 );
nor ( w3234 , w3233 , g5 );
nor ( w3235 , w3234 , g5 );
and ( w3236 , w4343 , g5 );
not ( w3237 , w3236 );
and ( w3238 , w3237 , g3 );
not ( w3239 , w3235 );
and ( w3240 , w3239 , w3238 );
nor ( w3241 , w3240 , g4 );
nor ( w3242 , w3241 , w1993 );
and ( w3243 , w3242 , g3 );
and ( w3244 , w3243 , w8728 );
nor ( w3245 , w3244 , w3072 );
nor ( w3246 , w3245 , g6 );
and ( w3247 , w3246 , w7997 );
and ( w3248 , w3247 , g2 );
and ( w3249 , w3248 , w8828 );
and ( w3250 , w3249 , w8765 );
and ( w3251 , w3250 , w8792 );
and ( w3252 , w8828 , g13 );
and ( w3253 , w3252 , w8845 );
and ( w3254 , w3251 , w3360 );
and ( w3255 , w3254 , w8837 );
nor ( w3256 , w3231 , w3255 );
not ( w3257 , w3256 );
and ( w3258 , w3257 , w400 );
not ( w3259 , w3258 );
and ( w3260 , w3259 , w3183 );
not ( w3261 , w3260 );
and ( w3262 , w3261 , g2 );
and ( w3263 , w8819 , w3197 );
and ( w3264 , w3263 , g10 );
and ( w3265 , w3264 , g12 );
and ( w3266 , w8819 , w3223 );
and ( w3267 , w3266 , g2 );
nor ( w3268 , w3265 , w3267 );
nor ( w3269 , w3268 , g16 );
and ( w3270 , w3269 , g15 );
and ( w3271 , w3270 , w400 );
and ( w3272 , w3271 , g14 );
not ( w3273 , w3272 );
and ( w3274 , w3273 , w3183 );
and ( w3275 , w5461 , w17 );
and ( w3276 , w3275 , w27 );
and ( w3277 , w3276 , g12 );
and ( w3278 , w3222 , w8828 );
and ( w3279 , w3278 , w7783 );
nor ( w3280 , w3277 , w3279 );
not ( w3281 , w3280 );
and ( w3282 , w3281 , g8 );
and ( w3283 , w3282 , g10 );
and ( w3284 , w2095 , w8735 );
and ( w3285 , w3284 , g10 );
and ( w3286 , w3285 , w8742 );
and ( w3287 , w3286 , g8 );
not ( w3288 , w3287 );
and ( w3289 , w3288 , w2190 );
and ( w3290 , w3289 , w7783 );
and ( w3291 , w3283 , w3290 );
nor ( w3292 , w3291 , g4 );
nor ( w3293 , w3292 , g13 );
and ( w3294 , w3200 , w8767 );
nor ( w3295 , w3294 , w566 );
nor ( w3296 , w3295 , g7 );
and ( w3297 , w3296 , w8769 );
and ( w3298 , w3297 , g10 );
and ( w3299 , w3298 , w33 );
and ( w3300 , w3299 , g12 );
and ( w3301 , w3222 , w7783 );
and ( w3302 , w3301 , w8837 );
nor ( w3303 , w3300 , w3302 );
not ( w3304 , w3303 );
and ( w3305 , w3304 , w2190 );
nor ( w3306 , w3305 , g4 );
nor ( w3307 , w3306 , g2 );
and ( w3308 , w3307 , w8819 );
and ( w3309 , w3308 , w8765 );
and ( w3310 , w3309 , w8845 );
and ( w3311 , w3310 , g15 );
and ( w3312 , w3311 , g14 );
and ( w3313 , w3312 , w8837 );
and ( w3314 , w3313 , w8828 );
nor ( w3315 , w3293 , w3314 );
nor ( w3316 , w3315 , g9 );
nor ( w3317 , w1578 , g10 );
not ( w3318 , w3317 );
and ( w3319 , w3318 , w1579 );
nor ( w3320 , w3319 , g8 );
nor ( w3321 , w3320 , g6 );
and ( w3322 , w3321 , g9 );
and ( w3323 , w3322 , w7783 );
and ( w3324 , w40 , w8767 );
and ( w3325 , w3324 , g9 );
and ( w3326 , w3325 , w1575 );
not ( w3327 , w3326 );
and ( w3328 , w3327 , g18 );
nor ( w3329 , w3328 , g6 );
and ( w3330 , w3329 , w1361 );
and ( w3331 , w3330 , w1579 );
nor ( w3332 , w3331 , g10 );
and ( w3333 , w3332 , w8767 );
nor ( w3334 , w3333 , g6 );
and ( w3335 , w3334 , w7783 );
and ( w3336 , w3323 , w3335 );
and ( w3337 , w3336 , w8792 );
nor ( w3338 , w3316 , w3337 );
nor ( w3339 , w3338 , g6 );
and ( w3340 , w3339 , g15 );
not ( w3341 , w3340 );
and ( w3342 , w3341 , w3183 );
nor ( w3343 , w3342 , g1 );
and ( w3344 , w3343 , w8828 );
and ( w3345 , w3344 , w7783 );
and ( w3346 , w3345 , g14 );
not ( w3347 , w3346 );
and ( w3348 , w3347 , w3183 );
nor ( w3349 , w3348 , g11 );
not ( w3350 , w3349 );
and ( w3351 , w3183 , w3350 );
and ( w3352 , w3274 , w3351 );
nor ( w3353 , w3352 , g11 );
nor ( w3354 , w3262 , w3353 );
nor ( w3355 , w3354 , g16 );
not ( w3356 , w3355 );
and ( w3357 , w3356 , w3183 );
nor ( w3358 , w3357 , g9 );
and ( w3359 , w3358 , w8792 );
not ( w3360 , w3253 );
and ( w3361 , w3359 , w3360 );
not ( w3362 , w3353 );
and ( w3363 , w3183 , w3362 );
not ( w3364 , w3361 );
and ( w3365 , w3364 , w3363 );
nor ( w3366 , w3365 , g11 );
not ( w3367 , w3366 );
and ( w3368 , w3183 , w3367 );
and ( w3369 , w7783 , w3368 );
and ( w3370 , w8767 , g6 );
and ( w3371 , w8845 , g9 );
nor ( w3372 , w2847 , w1423 );
and ( w3373 , w3372 , w408 );
nor ( w3374 , w3371 , w3373 );
not ( w3375 , w3374 );
and ( w3376 , w3375 , g2 );
and ( w3377 , w3376 , w8792 );
nor ( w3378 , w3370 , w3377 );
not ( w3379 , w3378 );
and ( w3380 , w3379 , g2 );
and ( w3381 , w3380 , w8792 );
and ( w3382 , w3381 , g11 );
not ( w3383 , w3382 );
and ( w3384 , w3115 , w3383 );
and ( w3385 , w3384 , g13 );
not ( w3386 , w3385 );
and ( w3387 , g13 , w3386 );
and ( w3388 , w3387 , g14 );
and ( w3389 , w3388 , g15 );
not ( w3390 , w3389 );
and ( w3391 , w3390 , w3115 );
and ( w3392 , w3391 , g16 );
and ( w3393 , w1 , g8 );
and ( w3394 , w3393 , w8735 );
and ( w3395 , w3394 , w8860 );
and ( w3396 , w3395 , w5461 );
nor ( w3397 , w3396 , g7 );
nor ( w3398 , w3397 , g5 );
and ( w3399 , w3398 , w17 );
and ( w3400 , w3399 , w8845 );
nor ( w3401 , w3400 , g5 );
not ( w3402 , w3401 );
and ( w3403 , w3402 , w27 );
nor ( w3404 , w3403 , g3 );
and ( w3405 , w3404 , w8860 );
nor ( w3406 , w3405 , g9 );
nor ( w3407 , w3406 , g9 );
nor ( w3408 , w15 , g7 );
nor ( w3409 , w3407 , w3408 );
and ( w3410 , w3409 , w8845 );
and ( w3411 , w3410 , g2 );
and ( w3412 , w3411 , w8792 );
nor ( w3413 , g6 , w3412 );
and ( w3414 , w3413 , g8 );
and ( w3415 , g13 , g6 );
nor ( w3416 , w3414 , w3415 );
and ( w3417 , w3416 , g10 );
and ( w3418 , w3417 , g14 );
and ( w3419 , w3418 , g15 );
not ( w3420 , w3419 );
and ( w3421 , w3420 , w3183 );
and ( w3422 , w3421 , w8828 );
not ( w3423 , w3422 );
and ( w3424 , w3423 , g10 );
and ( w3425 , w3424 , g2 );
and ( w3426 , w3425 , w8792 );
and ( w3427 , w3426 , g11 );
not ( w3428 , w3392 );
and ( w3429 , w3428 , w3427 );
and ( w3430 , w1354 , g14 );
and ( w3431 , w3430 , g15 );
and ( w3432 , w3431 , w8828 );
not ( w3433 , w3432 );
and ( w3434 , w3433 , w3183 );
and ( w3435 , w3183 , w3121 );
nor ( w3436 , w3435 , g10 );
and ( w3437 , w3436 , g15 );
not ( w3438 , w3437 );
and ( w3439 , w3438 , g15 );
and ( w3440 , w3439 , w8828 );
nor ( w3441 , w3434 , w3440 );
and ( w3442 , w3441 , g8 );
and ( w3443 , w8730 , g14 );
and ( w3444 , w3443 , g15 );
not ( w3445 , w3444 );
and ( w3446 , w3445 , w3115 );
and ( w3447 , w3446 , g16 );
nor ( w3448 , g6 , g13 );
and ( w3449 , w3677 , g17 );
nor ( w3450 , w3449 , g10 );
and ( w3451 , w7973 , w3450 );
and ( w3452 , w3451 , g11 );
nor ( w3453 , w3448 , w3452 );
and ( w3454 , w3453 , w3677 );
nor ( w3455 , w3454 , g10 );
and ( w3456 , w3455 , w8767 );
and ( w3457 , w3456 , g14 );
and ( w3458 , w3457 , g15 );
not ( w3459 , w3458 );
and ( w3460 , w3459 , w3183 );
and ( w3461 , w3460 , w8828 );
nor ( w3462 , w3461 , g10 );
and ( w3463 , w3462 , w8767 );
and ( w3464 , w3463 , g2 );
and ( w3465 , w3464 , w8792 );
and ( w3466 , w3465 , g11 );
not ( w3467 , w3447 );
and ( w3468 , w3467 , w3466 );
and ( w3469 , w1588 , w8767 );
and ( w3470 , w3469 , w8730 );
and ( w3471 , w3470 , w400 );
nor ( w3472 , w2844 , w3471 );
not ( w3473 , w3472 );
and ( w3474 , w3473 , w1361 );
not ( w3475 , w3474 );
and ( w3476 , w3475 , g13 );
and ( w3477 , w3476 , g16 );
nor ( w3478 , w3477 , g10 );
and ( w3479 , w3478 , w8767 );
and ( w3480 , w3479 , g2 );
and ( w3481 , w3480 , w8792 );
and ( w3482 , g13 , w3481 );
and ( w3483 , w3482 , g14 );
and ( w3484 , w3483 , g15 );
not ( w3485 , w3484 );
and ( w3486 , w3485 , w3115 );
and ( w3487 , w3486 , g16 );
and ( w3488 , w1414 , g14 );
and ( w3489 , w3488 , g15 );
and ( w3490 , w3489 , w8730 );
not ( w3491 , w3122 );
and ( w3492 , w3490 , w3491 );
not ( w3493 , w3121 );
and ( w3494 , w3492 , w3493 );
not ( w3495 , w3494 );
and ( w3496 , w3495 , w3183 );
and ( w3497 , w3496 , w8828 );
nor ( w3498 , w3497 , g8 );
and ( w3499 , w3498 , w8730 );
and ( w3500 , w3499 , w8792 );
not ( w3501 , w3487 );
and ( w3502 , w3501 , w3500 );
and ( w3503 , w3502 , g2 );
and ( w3504 , w3468 , w3503 );
nor ( w3505 , w3442 , w3504 );
nor ( w3506 , w3505 , g10 );
and ( w3507 , w3506 , g2 );
and ( w3508 , w3507 , g11 );
nor ( w3509 , w3429 , w3508 );
and ( w3510 , w519 , w8742 );
and ( w3511 , w3510 , w8769 );
and ( w3512 , w3511 , w8845 );
and ( w3513 , w3512 , w361 );
nor ( w3514 , w3513 , g7 );
and ( w3515 , w3514 , w8860 );
and ( w3516 , w3515 , w8769 );
and ( w3517 , w3516 , w8735 );
not ( w3518 , w3517 );
and ( w3519 , w3518 , w408 );
and ( w3520 , w3519 , g10 );
nor ( w3521 , w3520 , g9 );
nor ( w3522 , w3521 , g8 );
and ( w3523 , w3522 , w8845 );
nor ( w3524 , w3523 , g6 );
nor ( w3525 , w3524 , g1 );
and ( w3526 , w8860 , w59 );
and ( w3527 , w3526 , w3200 );
nor ( w3528 , w3527 , g5 );
nor ( w3529 , w3528 , g7 );
nor ( w3530 , w3529 , w270 );
not ( w3531 , w3530 );
and ( w3532 , w3531 , w361 );
nor ( w3533 , w3532 , g3 );
and ( w3534 , w3533 , w8765 );
and ( w3535 , w3534 , w8860 );
and ( w3536 , w1260 , w1220 );
nor ( w3537 , w3536 , g3 );
and ( w3538 , w3537 , w8765 );
nor ( w3539 , w3535 , w3538 );
and ( w3540 , w3539 , w8767 );
and ( w3541 , w361 , w1244 );
nor ( w3542 , w3541 , g9 );
and ( w3543 , w3542 , w8735 );
and ( w3544 , w3543 , w8860 );
not ( w3545 , w3544 );
and ( w3546 , w3545 , w1248 );
nor ( w3547 , w3546 , g5 );
and ( w3548 , w3547 , w8742 );
not ( w3549 , w3548 );
and ( w3550 , w3540 , w3549 );
and ( w3551 , w3550 , w8845 );
and ( w3552 , w3551 , w7783 );
and ( w3553 , w3552 , g10 );
nor ( w3554 , g6 , w3553 );
nor ( w3555 , w3554 , g2 );
and ( w3556 , w3525 , w3555 );
and ( w3557 , w3556 , g10 );
and ( w3558 , w3557 , w8767 );
and ( w3559 , w8792 , w1361 );
not ( w3560 , w3559 );
and ( w3561 , w3560 , g9 );
nor ( w3562 , w3561 , g1 );
and ( w3563 , g9 , w3562 );
and ( w3564 , w3563 , g6 );
not ( w3565 , w3564 );
and ( w3566 , w3565 , g6 );
nor ( w3567 , w3566 , g1 );
nor ( w3568 , g10 , g2 );
and ( w3569 , w3673 , g6 );
nor ( w3570 , w3569 , g8 );
and ( w3571 , w3570 , w8730 );
and ( w3572 , w3571 , w7783 );
and ( w3573 , w3567 , w3572 );
not ( w3574 , w3573 );
and ( w3575 , w3574 , g13 );
nor ( w3576 , w3575 , g2 );
not ( w3577 , w3576 );
and ( w3578 , w3577 , g16 );
nor ( w3579 , w3578 , g2 );
and ( w3580 , w3579 , w8792 );
nor ( w3581 , w3558 , w3580 );
nor ( w3582 , w3581 , g8 );
nor ( w3583 , g8 , w3582 );
nor ( w3584 , w3583 , g2 );
and ( w3585 , w3584 , w8792 );
and ( w3586 , g13 , w3585 );
not ( w3587 , w3586 );
and ( w3588 , w3587 , g16 );
not ( w3589 , w3588 );
and ( w3590 , w3589 , w40 );
and ( w3591 , w3590 , g14 );
and ( w3592 , w3591 , g15 );
not ( w3593 , w3592 );
and ( w3594 , w3593 , w3115 );
nor ( w3595 , w3594 , g1 );
and ( w3596 , w3595 , g11 );
not ( w3597 , w3596 );
and ( w3598 , w3597 , w3368 );
and ( w3599 , w3509 , w3598 );
and ( w3600 , w3599 , w8382 );
and ( w3601 , g17 , w8382 );
and ( w3602 , w8597 , w3368 );
and ( w3603 , w3602 , w3599 );
and ( w3604 , w3603 , g9 );
not ( w3605 , w3604 );
and ( w3606 , w3605 , g16 );
and ( w3607 , w3606 , w8833 );
and ( w3608 , w3607 , g1 );
not ( w3609 , w3608 );
and ( w3610 , w3609 , w3599 );
not ( w3611 , w3610 );
and ( w3612 , w3611 , g11 );
not ( w3613 , w3612 );
and ( w3614 , w3613 , w3368 );
nor ( w3615 , w3600 , w3614 );
and ( w3616 , w3615 , w8845 );
and ( w3617 , w3616 , w8833 );
and ( w3618 , w3617 , g1 );
not ( w3619 , w3618 );
and ( w3620 , w3619 , w3599 );
and ( w3621 , w3620 , g13 );
nor ( w3622 , w3621 , g15 );
and ( w3623 , w3622 , g1 );
not ( w3624 , w3623 );
and ( w3625 , w3624 , w3599 );
not ( w3626 , w3625 );
and ( w3627 , w3626 , g11 );
not ( w3628 , w3627 );
and ( w3629 , w3628 , w3368 );
nor ( w3630 , w3369 , w3629 );
and ( w3631 , w3630 , g13 );
not ( w3632 , w3631 );
and ( w3633 , w3632 , w3599 );
and ( w3634 , w17 , w8735 );
and ( w3635 , w3634 , w8860 );
and ( w3636 , w3635 , g10 );
and ( w3637 , w3636 , g12 );
and ( w3638 , w3637 , w8742 );
and ( w3639 , w3638 , w8837 );
and ( w3640 , w3639 , g8 );
and ( w3641 , w3640 , w8845 );
and ( w3642 , w3641 , w8819 );
and ( w3643 , w3585 , g11 );
and ( w3644 , w3643 , g13 );
nor ( w3645 , w3642 , w3644 );
not ( w3646 , w3645 );
and ( w3647 , w3646 , g15 );
and ( w3648 , w3647 , w7783 );
and ( w3649 , w3648 , g16 );
not ( w3650 , w3649 );
and ( w3651 , w3633 , w3650 );
not ( w3652 , w3651 );
and ( w3653 , w3652 , g14 );
nor ( w3654 , w3653 , w3084 );
and ( t_6 , w3654 , w3633 );
and ( w3655 , w2765 , w8860 );
and ( w3656 , w3655 , g10 );
and ( w3657 , w3656 , g12 );
and ( w3658 , w3657 , w8742 );
and ( w3659 , w3658 , w8837 );
and ( w3660 , w3659 , w8819 );
and ( w3661 , w3660 , g8 );
and ( w3662 , w3661 , g16 );
nor ( w3663 , w3662 , w1395 );
nor ( w3664 , w3663 , g6 );
and ( w3665 , w3664 , w8765 );
and ( w3666 , w3665 , g14 );
and ( w3667 , w3666 , w8168 );
not ( w3668 , w3667 );
and ( w3669 , w3668 , w1567 );
nor ( w3670 , w3669 , g1 );
and ( w3671 , w3670 , w7783 );
not ( w3672 , w3671 );
nand ( t_7 , w3672 , w1567 );
not ( w3673 , w3568 );
and ( w3674 , w3673 , w213 );
not ( w3675 , w3674 );
and ( w3676 , w3675 , g6 );
not ( w3677 , w2844 );
and ( w3678 , w40 , w3677 );
and ( w3679 , w3678 , w8730 );
nor ( w3680 , w3679 , g2 );
nor ( w3681 , w3680 , g10 );
and ( w3682 , w3681 , g11 );
nor ( w3683 , w2847 , w2669 );
nor ( w3684 , w3683 , g16 );
and ( w3685 , w3682 , w3684 );
and ( w3686 , w3685 , g14 );
and ( w3687 , w3686 , g15 );
and ( w3688 , w3687 , w8845 );
not ( w3689 , w3688 );
and ( w3690 , w3689 , g13 );
nor ( w3691 , w3690 , g16 );
nor ( w3692 , w3676 , w3691 );
and ( w3693 , w8374 , g10 );
not ( w3694 , w3693 );
and ( w3695 , w3694 , g2 );
and ( w3696 , w1515 , w7783 );
not ( w3697 , w3696 );
and ( w3698 , w3697 , g13 );
and ( w3699 , w3415 , w8828 );
and ( w3700 , w3699 , w33 );
and ( w3701 , w3700 , g15 );
and ( w3702 , w3701 , g14 );
and ( w3703 , g4 , w8819 );
and ( w3704 , w3703 , w8735 );
and ( w3705 , w3704 , w8837 );
and ( w3706 , w3705 , w7997 );
and ( w3707 , w3706 , w8828 );
and ( w3708 , w3707 , w8765 );
and ( w3709 , w3448 , g2 );
nor ( w3710 , g3 , g13 );
and ( w3711 , w3710 , w7783 );
and ( w3712 , w3711 , w8837 );
and ( w3713 , w3712 , w8828 );
and ( w3714 , w3713 , w8765 );
and ( w3715 , w3714 , w7141 );
and ( w3716 , w3714 , w122 );
and ( w3717 , w3716 , g12 );
and ( w3718 , w3717 , w8860 );
nor ( w3719 , w3715 , w3718 );
not ( w3720 , w3719 );
and ( w3721 , w3720 , g12 );
and ( w3722 , w3721 , w8860 );
nor ( w3723 , w3709 , w3722 );
and ( w3724 , w3723 , w8860 );
not ( w3725 , w3724 );
and ( w3726 , w3725 , g12 );
and ( w3727 , w3726 , w8837 );
and ( w3728 , w3727 , w7997 );
and ( w3729 , w3728 , w8828 );
and ( w3730 , w3729 , w8765 );
and ( w3731 , w3730 , w8845 );
and ( w3732 , w3731 , w8735 );
and ( w3733 , w3732 , w8819 );
and ( w3734 , w3733 , g2 );
not ( w3735 , w1846 );
and ( w3736 , w3735 , g4 );
and ( w3737 , w3736 , w8837 );
and ( w3738 , w3737 , w8728 );
and ( w3739 , w3730 , w8735 );
and ( w3740 , w3739 , g4 );
nor ( w3741 , w3740 , w3722 );
nor ( w3742 , w3741 , g13 );
and ( w3743 , w3742 , w7783 );
nor ( w3744 , w3738 , w3743 );
nor ( w3745 , w3744 , g13 );
and ( w3746 , w3745 , w7997 );
and ( w3747 , w3746 , w8828 );
and ( w3748 , w3747 , w8765 );
and ( w3749 , w3748 , w8845 );
nor ( w3750 , w3722 , w3749 );
not ( w3751 , w3734 );
and ( w3752 , w3751 , w3750 );
not ( w3753 , w3058 );
and ( w3754 , w3753 , w3752 );
nor ( w3755 , w3754 , g13 );
and ( w3756 , w3755 , w8860 );
and ( w3757 , w3756 , g2 );
not ( w3758 , w3757 );
and ( w3759 , w3758 , w3750 );
nor ( w3760 , w3759 , g11 );
and ( w3761 , w3760 , w7997 );
and ( w3762 , w3761 , w8828 );
nor ( w3763 , w3708 , w3762 );
not ( w3764 , w3763 );
and ( w3765 , w3764 , g2 );
not ( w3766 , w3765 );
and ( w3767 , w3766 , w3750 );
nor ( w3768 , w122 , g7 );
not ( w3769 , w3768 );
and ( w3770 , w3769 , g11 );
and ( w3771 , w3770 , w7997 );
not ( w3772 , w3771 );
and ( w3773 , w3772 , w3767 );
not ( w3774 , w3773 );
and ( w3775 , w3774 , g6 );
and ( w3776 , w3775 , w8819 );
and ( w3777 , w3776 , w8765 );
and ( w3778 , w3777 , w8828 );
not ( w3779 , w3778 );
and ( w3780 , w3767 , w3779 );
not ( w3781 , w3780 );
and ( w3782 , w3781 , g2 );
and ( w3783 , w289 , g8 );
and ( w3784 , w3783 , w8742 );
and ( w3785 , w3784 , w59 );
nor ( w3786 , w3785 , g5 );
not ( w3787 , w3786 );
and ( w3788 , w3787 , g10 );
and ( w3789 , w3788 , w8742 );
nor ( w3790 , w3789 , g7 );
not ( w3791 , w3790 );
and ( w3792 , w3791 , w13 );
not ( w3793 , w3792 );
and ( w3794 , w3793 , g8 );
nor ( w3795 , w79 , w3794 );
and ( w3796 , w3795 , w8735 );
and ( w3797 , w3796 , w8860 );
and ( w3798 , w3797 , g2 );
and ( w3799 , w3798 , w2585 );
and ( w3800 , w8735 , g11 );
and ( w3801 , w514 , w8860 );
and ( w3802 , w3801 , w8728 );
and ( w3803 , w3802 , w8765 );
and ( w3804 , w3803 , w8819 );
and ( w3805 , w3804 , w8828 );
and ( w3806 , w516 , w8828 );
and ( w3807 , w3806 , w8728 );
and ( w3808 , w3807 , g13 );
and ( w3809 , w3808 , g11 );
not ( w3810 , w3809 );
and ( w3811 , w3810 , w3767 );
nor ( w3812 , w3811 , w213 );
nor ( w3813 , w3805 , w3812 );
nor ( w3814 , w3813 , g3 );
and ( w3815 , w3814 , g11 );
not ( w3816 , w3815 );
and ( w3817 , w3816 , w3767 );
nor ( w3818 , w3817 , w213 );
nor ( w3819 , w3800 , w3818 );
nor ( w3820 , w3819 , g4 );
and ( w3821 , w3820 , g6 );
nor ( w3822 , w3821 , w3818 );
nor ( w3823 , w3822 , g13 );
nor ( w3824 , w3823 , w3812 );
nor ( w3825 , w3824 , g3 );
and ( w3826 , w3825 , w8765 );
and ( w3827 , w3826 , w8828 );
and ( w3828 , w3827 , w8728 );
and ( w3829 , w3828 , w7783 );
and ( w3830 , w3829 , g11 );
and ( w3831 , w551 , w8168 );
nor ( w3832 , w3831 , g7 );
nor ( w3833 , w3832 , g7 );
and ( w3834 , w3833 , w7141 );
not ( w3835 , w3834 );
and ( w3836 , w3835 , g11 );
nor ( w3837 , w3836 , w3818 );
not ( w3838 , w3837 );
and ( w3839 , w3838 , g2 );
and ( w3840 , w3827 , g14 );
and ( w3841 , w3840 , w7783 );
and ( w3842 , w3841 , g6 );
nor ( w3843 , w3842 , w3818 );
not ( w3844 , w3839 );
and ( w3845 , w3844 , w3843 );
nor ( w3846 , w3845 , g10 );
and ( w3847 , w3846 , g6 );
nor ( w3848 , w3847 , w3818 );
nor ( w3849 , w3848 , g13 );
nor ( w3850 , w3849 , w3812 );
nor ( w3851 , w3850 , g3 );
and ( w3852 , w3851 , w8765 );
and ( w3853 , w3852 , w8828 );
not ( w3854 , w3853 );
and ( w3855 , w3767 , w3854 );
not ( w3856 , w3830 );
and ( w3857 , w3856 , w3855 );
not ( w3858 , w3857 );
and ( w3859 , w3858 , g10 );
nor ( w3860 , w3859 , w3853 );
not ( w3861 , w3860 );
and ( w3862 , w3861 , g6 );
nor ( w3863 , w3862 , w3818 );
nor ( w3864 , w3863 , g3 );
nor ( w3865 , w3799 , w3864 );
not ( w3866 , w3865 );
and ( w3867 , w3866 , w779 );
and ( w3868 , w3867 , g6 );
and ( w3869 , w3868 , g11 );
not ( w3870 , w3869 );
and ( w3871 , w3870 , w3855 );
not ( w3872 , w3871 );
and ( w3873 , w3872 , w33 );
nor ( w3874 , w3873 , w3853 );
not ( w3875 , w3874 );
and ( w3876 , w3875 , g6 );
nor ( w3877 , w3876 , w3818 );
nor ( w3878 , w3877 , g13 );
nor ( w3879 , w3878 , w3812 );
nor ( w3880 , w3879 , g3 );
and ( w3881 , w3880 , w8765 );
and ( w3882 , w3881 , w8828 );
nor ( w3883 , g4 , w3882 );
not ( w3884 , w3883 );
and ( w3885 , w3884 , g11 );
not ( w3886 , w3885 );
and ( w3887 , w3886 , w3855 );
not ( w3888 , w3887 );
and ( w3889 , w3888 , g10 );
nor ( w3890 , w3889 , w3853 );
not ( w3891 , w3890 );
and ( w3892 , w3891 , g6 );
nor ( w3893 , w3892 , w3818 );
nor ( w3894 , w3893 , g13 );
nor ( w3895 , w3894 , w3812 );
nor ( w3896 , w3895 , g3 );
and ( w3897 , w3896 , w8765 );
and ( w3898 , w3897 , w8828 );
not ( w3899 , w3898 );
and ( w3900 , w3899 , w3767 );
not ( w3901 , w3782 );
and ( w3902 , w3901 , w3900 );
nor ( w3903 , w3902 , g3 );
and ( w3904 , w3903 , w8728 );
not ( w3905 , w3904 );
and ( w3906 , w3905 , w3900 );
and ( w3907 , w3906 , g13 );
and ( w3908 , w3994 , g14 );
and ( w3909 , w3908 , g15 );
nor ( w3910 , w299 , w1244 );
not ( w3911 , w3910 );
and ( w3912 , w3911 , g3 );
and ( w3913 , w3912 , w8765 );
and ( w3914 , w3913 , w8828 );
nor ( w3915 , g4 , w3914 );
not ( w3916 , w3915 );
and ( w3917 , w3916 , g3 );
and ( w3918 , w3917 , w8765 );
and ( w3919 , w3918 , w8828 );
and ( w3920 , w473 , g2 );
nor ( w3921 , g11 , g2 );
and ( w3922 , w3921 , w8819 );
nor ( w3923 , w3920 , w3922 );
not ( w3924 , w245 );
and ( w3925 , w3924 , g2 );
not ( w3926 , w244 );
and ( w3927 , w3926 , g2 );
nor ( w3928 , w3927 , g6 );
and ( w3929 , w3928 , w8735 );
and ( w3930 , w3929 , w8765 );
not ( w3931 , w3925 );
and ( w3932 , w3931 , w3930 );
and ( w3933 , w3932 , g8 );
not ( w3934 , w3933 );
and ( w3935 , w3934 , g8 );
not ( w3936 , w3935 );
and ( w3937 , w3936 , w779 );
and ( w3938 , w3937 , w8735 );
and ( w3939 , w3938 , w8765 );
not ( w3940 , w3923 );
and ( w3941 , w3940 , w3939 );
and ( w3942 , w3941 , w8769 );
and ( w3943 , w3942 , w8845 );
and ( w3944 , w3943 , w8742 );
and ( w3945 , w3944 , g8 );
and ( w3946 , w1609 , g12 );
and ( w3947 , w3946 , w8742 );
and ( w3948 , w3947 , g8 );
not ( w3949 , w3945 );
and ( w3950 , w3949 , w3948 );
not ( w3951 , w3950 );
and ( w3952 , w3951 , w770 );
and ( w3953 , w3952 , w8819 );
and ( w3954 , w3953 , w8742 );
and ( w3955 , w3954 , g10 );
and ( w3956 , w3955 , w8769 );
and ( w3957 , w3956 , g14 );
and ( w3958 , w3957 , w779 );
and ( w3959 , w3958 , w33 );
and ( w3960 , w3959 , w17 );
and ( w3961 , w3960 , w8828 );
nor ( w3962 , w3961 , w3699 );
not ( w3963 , w3962 );
and ( w3964 , w3963 , g10 );
and ( w3965 , w3964 , w8769 );
and ( w3966 , w3965 , g14 );
and ( w3967 , w3966 , w33 );
and ( w3968 , w3967 , w59 );
and ( w3969 , w3968 , w8860 );
and ( w3970 , w3969 , w8735 );
and ( w3971 , w3970 , w8765 );
nor ( w3972 , w3971 , g5 );
and ( w3973 , w3972 , w8742 );
and ( w3974 , w3973 , w8860 );
and ( w3975 , w3971 , w8845 );
not ( w3976 , w3975 );
and ( w3977 , w3976 , w3948 );
and ( w3978 , w3971 , w8767 );
nor ( w3979 , w3978 , g8 );
nor ( w3980 , w3979 , g7 );
and ( w3981 , w3980 , g14 );
and ( w3982 , w3981 , w33 );
and ( w3983 , w3982 , w17 );
and ( w3984 , w3983 , w27 );
and ( w3985 , w3984 , w8828 );
not ( w3986 , w3977 );
and ( w3987 , w3986 , w3985 );
nor ( w3988 , w3987 , w3699 );
not ( w3989 , w3988 );
and ( w3990 , w3989 , g14 );
and ( w3991 , w3990 , g15 );
and ( w3992 , w3991 , w33 );
and ( w3993 , w3992 , g12 );
not ( w3994 , w3907 );
and ( w3995 , w3994 , w3993 );
nor ( w3996 , g7 , w1786 );
nor ( w3997 , w3996 , g3 );
and ( w3998 , w3997 , w8765 );
and ( w3999 , w3998 , w33 );
and ( w4000 , w92 , w8845 );
and ( w4001 , w4000 , w8819 );
and ( w4002 , w4001 , w8828 );
nor ( w4003 , w3999 , w4002 );
and ( w4004 , w4003 , w213 );
nor ( w4005 , w121 , w4002 );
nor ( w4006 , w4005 , g16 );
not ( w4007 , w4004 );
and ( w4008 , w4007 , w4006 );
and ( w4009 , w4008 , w8845 );
and ( w4010 , w4009 , w8819 );
not ( w4011 , w4010 );
and ( w4012 , w4011 , w3906 );
not ( w4013 , w4012 );
and ( w4014 , w4013 , g2 );
and ( w4015 , w4014 , g11 );
nor ( w4016 , w1395 , g10 );
nor ( w4017 , w4016 , g10 );
not ( w4018 , w4017 );
and ( w4019 , w4018 , g15 );
not ( w4020 , w4019 );
and ( w4021 , w4020 , g15 );
not ( w4022 , w4021 );
and ( w4023 , w4022 , g7 );
and ( w4024 , w1786 , w8819 );
nor ( w4025 , w4024 , w3699 );
not ( w4026 , w4025 );
and ( w4027 , w4026 , g5 );
and ( w4028 , w4027 , w33 );
nor ( w4029 , w4028 , w4002 );
not ( w4030 , w4029 );
and ( w4031 , w4030 , g14 );
and ( w4032 , w4031 , g15 );
and ( w4033 , w4032 , g12 );
and ( w4034 , w4033 , w8735 );
and ( w4035 , w4034 , w8765 );
and ( w4036 , w4035 , w8828 );
and ( w4037 , w4036 , g2 );
nor ( w4038 , w4023 , w4037 );
nor ( w4039 , w4038 , g13 );
and ( w4040 , w4039 , g14 );
and ( w4041 , w4040 , g2 );
and ( w4042 , w4041 , w8837 );
not ( w4043 , w4042 );
and ( w4044 , w4043 , w3767 );
not ( w4045 , w4044 );
and ( w4046 , w4045 , g2 );
and ( w4047 , w4046 , g12 );
and ( w4048 , w4047 , w8735 );
and ( w4049 , w4048 , w8765 );
and ( w4050 , w4049 , w8828 );
nor ( w4051 , w4015 , w4050 );
nor ( w4052 , w3997 , w92 );
and ( w4053 , w4052 , w213 );
nor ( w4054 , w4053 , g3 );
and ( w4055 , w4054 , w8845 );
and ( w4056 , w4055 , g11 );
not ( w4057 , w3714 );
and ( w4058 , w4057 , w3767 );
nor ( w4059 , w4058 , g10 );
and ( w4060 , w4059 , w7783 );
and ( w4061 , w4060 , w8735 );
nor ( w4062 , w1786 , w4061 );
nor ( w4063 , w4062 , g6 );
and ( w4064 , w4063 , g14 );
and ( w4065 , w4064 , w8837 );
not ( w4066 , w4065 );
and ( w4067 , w4066 , w3767 );
nor ( w4068 , w4067 , g2 );
and ( w4069 , w4068 , g12 );
and ( w4070 , w4069 , w8765 );
and ( w4071 , w4070 , w8828 );
not ( w4072 , w4071 );
and ( w4073 , w4072 , w3767 );
and ( w4074 , w5920 , w4073 );
nor ( w4075 , w4074 , g11 );
and ( w4076 , w4075 , w7783 );
and ( w4077 , w4076 , g12 );
and ( w4078 , w4077 , w8765 );
and ( w4079 , w4078 , w8828 );
nor ( w4080 , w4056 , w4079 );
nor ( w4081 , w4080 , g13 );
and ( w4082 , w4081 , w7783 );
and ( w4083 , w4082 , g12 );
and ( w4084 , w4083 , w8860 );
and ( w4085 , w4084 , w8765 );
and ( w4086 , w4085 , w8828 );
not ( w4087 , w4086 );
and ( w4088 , w4051 , w4087 );
not ( w4089 , w4088 );
and ( w4090 , w4089 , g12 );
and ( w4091 , w4090 , w27 );
not ( w4092 , w4091 );
and ( w4093 , w4092 , w3906 );
nor ( w4094 , w4093 , g3 );
and ( w4095 , w4094 , w8765 );
nor ( w4096 , w3995 , w4095 );
and ( w4097 , w4096 , w3906 );
and ( w4098 , w8860 , w4097 );
and ( w4099 , w8769 , g12 );
and ( w4100 , w4099 , w8742 );
and ( w4101 , w4098 , w4110 );
not ( w4102 , w4101 );
and ( w4103 , w4102 , g7 );
nor ( w4104 , w4100 , w4037 );
not ( w4105 , w4104 );
and ( w4106 , w4105 , g5 );
nor ( w4107 , w4106 , w3971 );
and ( w4108 , w4107 , w8860 );
and ( w4109 , w4108 , g2 );
not ( w4110 , w4100 );
and ( w4111 , w4097 , w4110 );
and ( w4112 , w4111 , g2 );
not ( w4113 , w4112 );
and ( w4114 , w4113 , w1786 );
nor ( w4115 , w4114 , w3971 );
and ( w4116 , w4115 , g12 );
and ( w4117 , w4116 , w4245 );
and ( w4118 , w3992 , w27 );
not ( w4119 , w4118 );
and ( w4120 , g10 , w4119 );
and ( w4121 , w4120 , w8860 );
and ( w4122 , w4121 , w8769 );
and ( w4123 , w4122 , w8742 );
and ( w4124 , w4123 , w3767 );
nor ( w4125 , w4117 , w4124 );
and ( w4126 , w4125 , g14 );
and ( w4127 , w4126 , g15 );
not ( w4128 , w1260 );
and ( w4129 , w4128 , w4097 );
not ( w4130 , w4129 );
and ( w4131 , w4130 , w299 );
and ( w4132 , w4006 , w8742 );
nor ( w4133 , w4131 , w4132 );
nor ( w4134 , w4133 , g3 );
not ( w4135 , w4134 );
and ( w4136 , w4135 , g12 );
not ( w4137 , w4136 );
and ( w4138 , w4137 , g5 );
and ( w4139 , w4138 , w8845 );
and ( w4140 , w4139 , w8735 );
and ( w4141 , w4140 , w8819 );
not ( w4142 , w4141 );
and ( w4143 , w4142 , w3906 );
nor ( w4144 , w4143 , g3 );
and ( w4145 , w4144 , w8765 );
and ( w4146 , w4145 , w8828 );
not ( w4147 , w4146 );
and ( w4148 , w3120 , w4147 );
and ( w4149 , w1898 , w3200 );
not ( w4150 , w4148 );
and ( w4151 , w4150 , w4149 );
not ( w4152 , w4151 );
and ( w4153 , w4152 , w4097 );
not ( w4154 , w4153 );
and ( w4155 , w4154 , w299 );
nor ( w4156 , w4155 , w4132 );
nor ( w4157 , w4156 , g3 );
not ( w4158 , w4157 );
and ( w4159 , w4158 , g12 );
nor ( w4160 , w4159 , g3 );
and ( w4161 , w4160 , g5 );
nor ( w4162 , g4 , w122 );
and ( w4163 , w4162 , g2 );
and ( w4164 , w4163 , w7141 );
nor ( w4165 , w224 , w122 );
nor ( w4166 , g3 , w4165 );
and ( w4167 , w4166 , w8860 );
nor ( w4168 , w4167 , g4 );
not ( w4169 , w4168 );
and ( w4170 , w4169 , w400 );
nor ( w4171 , w4170 , w1260 );
and ( w4172 , g7 , g2 );
and ( w4173 , w4172 , w8730 );
not ( w4174 , w4173 );
and ( w4175 , w4174 , g2 );
not ( w4176 , w4175 );
and ( w4177 , w4176 , g15 );
and ( w4178 , w4177 , w1609 );
not ( w4179 , w4178 );
and ( w4180 , w4179 , g15 );
and ( w4181 , w4180 , w8860 );
nor ( w4182 , w4171 , w4181 );
and ( w4183 , w4182 , w8845 );
nor ( w4184 , g3 , g7 );
nor ( w4185 , w4183 , w4184 );
nor ( w4186 , w4185 , g3 );
and ( w4187 , w4186 , w8769 );
and ( w4188 , w4187 , w8845 );
not ( w4189 , w4164 );
and ( w4190 , w4189 , w4188 );
nor ( w4191 , w4190 , w4184 );
and ( w4192 , w4191 , w8728 );
nor ( w4193 , w4192 , g3 );
and ( w4194 , w4193 , w8769 );
and ( w4195 , w4194 , w8730 );
and ( w4196 , w4195 , w8845 );
and ( w4197 , w4196 , w8828 );
nor ( w4198 , w4161 , w4197 );
nor ( w4199 , w4198 , g10 );
and ( w4200 , w4199 , w8845 );
and ( w4201 , w4200 , w8819 );
not ( w4202 , w4201 );
and ( w4203 , w4202 , w3906 );
nor ( w4204 , w4203 , g3 );
and ( w4205 , w4204 , w408 );
not ( w4206 , w4205 );
and ( w4207 , w4206 , w3906 );
not ( w4208 , w4207 );
and ( w4209 , w4208 , w361 );
and ( w4210 , w4209 , w8828 );
nor ( w4211 , w121 , w4210 );
nor ( w4212 , w4211 , g6 );
and ( w4213 , w4212 , g11 );
and ( w4214 , w4213 , w7997 );
not ( w4215 , w4214 );
and ( w4216 , w4215 , w3767 );
nor ( w4217 , w4216 , g13 );
not ( w4218 , w4217 );
and ( w4219 , w4218 , w3906 );
nor ( w4220 , w4219 , g3 );
and ( w4221 , w4220 , w8765 );
and ( w4222 , w4221 , w8828 );
nor ( w4223 , w4127 , w4222 );
nor ( w4224 , w4223 , g13 );
not ( w4225 , w4224 );
and ( w4226 , w4225 , w3906 );
nor ( w4227 , w4226 , g3 );
and ( w4228 , w4227 , w8765 );
and ( w4229 , w4228 , w8828 );
nor ( w4230 , g4 , w4229 );
nor ( w4231 , w4230 , w4124 );
and ( w4232 , w4231 , g14 );
and ( w4233 , w4232 , g15 );
nor ( w4234 , w4233 , w4222 );
nor ( w4235 , w4234 , g13 );
not ( w4236 , w4235 );
and ( w4237 , w4236 , w3906 );
nor ( w4238 , w4237 , g3 );
and ( w4239 , w4238 , w8765 );
and ( w4240 , w4239 , w8828 );
not ( w4241 , w4109 );
and ( w4242 , w4241 , w4240 );
not ( w4243 , w4242 );
and ( w4244 , w4243 , g12 );
not ( w4245 , w4002 );
and ( w4246 , w4244 , w4245 );
nor ( w4247 , w4246 , w4124 );
and ( w4248 , w4247 , g14 );
and ( w4249 , w4248 , g15 );
nor ( w4250 , w4249 , w4222 );
nor ( w4251 , w4250 , g13 );
not ( w4252 , w4251 );
and ( w4253 , w4252 , w3906 );
nor ( w4254 , w4253 , g3 );
and ( w4255 , w4254 , w8765 );
and ( w4256 , w4255 , w8828 );
nor ( w4257 , w4103 , w4256 );
and ( w4258 , w4257 , g12 );
nor ( w4259 , w4258 , w4124 );
and ( w4260 , w4259 , g14 );
and ( w4261 , w4260 , g15 );
nor ( w4262 , w4261 , w4222 );
nor ( w4263 , w4262 , g13 );
not ( w4264 , w4263 );
and ( w4265 , w4264 , w3906 );
nor ( w4266 , w4265 , g3 );
and ( w4267 , w4266 , w8765 );
and ( w4268 , w4267 , w8828 );
not ( w4269 , w3974 );
and ( w4270 , w4269 , w4268 );
nor ( w4271 , w4118 , g5 );
and ( w4272 , w4271 , w8860 );
and ( w4273 , w4272 , w8742 );
and ( w4274 , w4273 , w3767 );
not ( w4275 , w4274 );
and ( w4276 , w4270 , w4275 );
nor ( w4277 , w4276 , w4002 );
not ( w4278 , w4277 );
and ( w4279 , w4278 , g14 );
and ( w4280 , w4279 , g15 );
nor ( w4281 , w4280 , w4222 );
nor ( w4282 , w4281 , g9 );
and ( w4283 , w4282 , w8819 );
not ( w4284 , w4283 );
and ( w4285 , w4284 , w3906 );
not ( w4286 , w3919 );
and ( w4287 , w4286 , w4285 );
nor ( w4288 , w4287 , g13 );
not ( w4289 , w4288 );
and ( w4290 , w4289 , w4285 );
nor ( w4291 , w4290 , w213 );
and ( w4292 , w4291 , g6 );
and ( w4293 , w3448 , w7997 );
and ( w4294 , w4293 , w8828 );
nor ( w4295 , w3909 , w4294 );
nor ( w4296 , w4295 , g6 );
and ( w4297 , w4296 , g11 );
and ( w4298 , w4297 , g3 );
not ( w4299 , w4298 );
and ( w4300 , w4299 , w4285 );
nor ( w4301 , w4300 , g9 );
and ( w4302 , w4301 , w8828 );
nor ( w4303 , w4292 , w4302 );
not ( w4304 , w4303 );
and ( w4305 , w4304 , g11 );
not ( w4306 , w4305 );
and ( w4307 , w4306 , w4285 );
and ( w4308 , g11 , w8742 );
and ( w4309 , w4308 , w8860 );
and ( w4310 , w4309 , w8769 );
and ( w4311 , w4310 , g6 );
and ( w4312 , w4311 , w8819 );
and ( w4313 , w4312 , w7997 );
not ( w4314 , w4313 );
and ( w4315 , w4314 , w3767 );
nor ( w4316 , w4315 , g1 );
and ( w4317 , w4316 , w8765 );
and ( w4318 , w4317 , w8828 );
and ( w4319 , w4307 , w4691 );
not ( w4320 , w4319 );
and ( w4321 , w4320 , g2 );
not ( w4322 , w162 );
and ( w4323 , w4322 , w4285 );
nor ( w4324 , w4323 , g6 );
and ( w4325 , w4324 , g3 );
not ( w4326 , w4325 );
and ( w4327 , w4326 , w4285 );
nor ( w4328 , w4327 , g9 );
and ( w4329 , w4328 , w8828 );
and ( w4330 , w4329 , g14 );
and ( w4331 , w4330 , g15 );
and ( w4332 , w4331 , g3 );
not ( w4333 , w4332 );
and ( w4334 , w4333 , w4285 );
and ( w4335 , w4334 , w8845 );
nor ( w4336 , w381 , g6 );
and ( w4337 , w4336 , g13 );
nor ( w4338 , w4337 , g16 );
not ( w4339 , w4335 );
and ( w4340 , w4339 , w4338 );
and ( w4341 , w4340 , g14 );
and ( w4342 , w4341 , g15 );
not ( w4343 , w476 );
and ( w4344 , w4343 , w4285 );
nor ( w4345 , w4344 , w213 );
and ( w4346 , w4345 , w4338 );
and ( w4347 , w4346 , w8845 );
and ( w4348 , w4347 , g11 );
nor ( w4349 , w4348 , g12 );
nor ( w4350 , w204 , g10 );
not ( w4351 , w4350 );
and ( w4352 , w4351 , g2 );
and ( w4353 , w4352 , w8845 );
and ( w4354 , w4353 , g11 );
not ( w4355 , w4354 );
and ( w4356 , w4355 , w4285 );
and ( w4357 , g10 , g6 );
not ( w4358 , w40 );
and ( w4359 , w4358 , g2 );
and ( w4360 , w4359 , w8845 );
and ( w4361 , w4360 , w400 );
and ( w4362 , w4361 , w8845 );
nor ( w4363 , w4362 , g6 );
nor ( w4364 , w4363 , g10 );
nor ( w4365 , w4364 , g10 );
not ( w4366 , w4365 );
and ( w4367 , w4366 , g11 );
nor ( w4368 , w4367 , g2 );
and ( w4369 , w4368 , g3 );
and ( w4370 , w4369 , g14 );
and ( w4371 , w4370 , g15 );
not ( w4372 , w4371 );
and ( w4373 , w4372 , w4285 );
nor ( w4374 , w4373 , g9 );
and ( w4375 , w4374 , w8828 );
nor ( w4376 , w4357 , w4375 );
and ( w4377 , w4376 , g11 );
and ( w4378 , w2844 , w8837 );
nor ( w4379 , w4377 , w4378 );
and ( w4380 , w4379 , w3684 );
and ( w4381 , w4380 , w8792 );
not ( w4382 , w4381 );
and ( w4383 , w4382 , g13 );
not ( w4384 , w4383 );
and ( w4385 , w4384 , g14 );
and ( w4386 , w4385 , g15 );
and ( w4387 , w4386 , g3 );
not ( w4388 , w4387 );
and ( w4389 , w4388 , w4285 );
nor ( w4390 , w4389 , g16 );
and ( w4391 , w4390 , w7783 );
and ( w4392 , w4391 , w3684 );
not ( w4393 , w4392 );
and ( w4394 , w4393 , g13 );
not ( w4395 , w4394 );
and ( w4396 , w4395 , g14 );
and ( w4397 , w4396 , g15 );
and ( w4398 , w4397 , g3 );
not ( w4399 , w4398 );
and ( w4400 , w4399 , w4285 );
nor ( w4401 , w4400 , g9 );
and ( w4402 , w4401 , w8828 );
not ( w4403 , w4402 );
and ( w4404 , w4356 , w4403 );
and ( w4405 , w4404 , g13 );
not ( w4406 , w4405 );
and ( w4407 , w4406 , g14 );
and ( w4408 , w4407 , g15 );
and ( w4409 , w4408 , g3 );
not ( w4410 , w4409 );
and ( w4411 , w4410 , w4285 );
nor ( w4412 , w4411 , g16 );
and ( w4413 , w4412 , w8765 );
and ( w4414 , w4413 , g14 );
and ( w4415 , w4414 , g15 );
and ( w4416 , w1516 , w8765 );
and ( w4417 , w4416 , w8730 );
and ( w4418 , w8730 , g4 );
and ( w4419 , w4418 , w7783 );
and ( w4420 , w4417 , w4419 );
not ( w4421 , w4420 );
and ( w4422 , w4421 , w4285 );
not ( w4423 , w4422 );
and ( w4424 , w4423 , g6 );
not ( w4425 , w4424 );
and ( w4426 , w4425 , g13 );
not ( w4427 , w4426 );
and ( w4428 , w4427 , g4 );
and ( w4429 , w4428 , g3 );
and ( w4430 , w4429 , g11 );
and ( w4431 , w4430 , w7997 );
not ( w4432 , w4431 );
and ( w4433 , w4432 , w3767 );
not ( w4434 , w4433 );
and ( w4435 , w4434 , g3 );
and ( w4436 , w4435 , w408 );
not ( w4437 , w4436 );
and ( w4438 , w4437 , w4285 );
nor ( w4439 , w4438 , g16 );
and ( w4440 , g4 , w4439 );
and ( w4441 , w4285 , w7783 );
and ( w4442 , w4441 , g13 );
and ( w4443 , g2 , g13 );
nor ( w4444 , w4443 , g16 );
and ( w4445 , w4444 , g6 );
nor ( w4446 , w4445 , w4294 );
and ( w4447 , w4446 , g14 );
not ( w4448 , w2619 );
and ( w4449 , w4448 , g6 );
and ( w4450 , w5243 , g6 );
nor ( w4451 , w4450 , w4294 );
nor ( w4452 , w4451 , g1 );
and ( w4453 , w4452 , w7997 );
and ( w4454 , w4453 , w8765 );
and ( w4455 , w4454 , w8828 );
not ( w4456 , w4447 );
and ( w4457 , w4456 , w4455 );
and ( w4458 , w4457 , g3 );
and ( w4459 , w4458 , g11 );
not ( w4460 , w4459 );
and ( w4461 , w4460 , w3767 );
and ( w4462 , w4461 , g12 );
not ( w4463 , w4462 );
and ( w4464 , w4463 , g3 );
not ( w4465 , w4464 );
and ( w4466 , w4465 , w4285 );
nor ( w4467 , w4466 , g9 );
and ( w4468 , w4467 , w8828 );
not ( w4469 , w4442 );
and ( w4470 , w4469 , w4468 );
nor ( w4471 , w4470 , g15 );
and ( w4472 , g10 , w8742 );
not ( w4473 , w4472 );
and ( w4474 , w4473 , g10 );
and ( w4475 , w2619 , g3 );
and ( w4476 , w4475 , w8792 );
and ( w4477 , w2077 , w3767 );
not ( w4478 , w4477 );
and ( w4479 , w4478 , g3 );
and ( w4480 , w4479 , w408 );
not ( w4481 , w4480 );
and ( w4482 , w4481 , w4285 );
not ( w4483 , w4482 );
and ( w4484 , w4476 , w4483 );
not ( w4485 , w4484 );
and ( w4486 , w4485 , g13 );
and ( w4487 , w4486 , w8168 );
nor ( w4488 , w4487 , w213 );
and ( w4489 , w4488 , g3 );
not ( w4490 , w4489 );
and ( w4491 , w4490 , w4285 );
nor ( w4492 , w4491 , g9 );
and ( w4493 , w4492 , w8828 );
not ( w4494 , w4474 );
and ( w4495 , w4494 , w4493 );
and ( w4496 , w4495 , w8792 );
and ( w4497 , w4496 , w8860 );
and ( w4498 , w4497 , g6 );
and ( w4499 , w4498 , w1489 );
nor ( w4500 , w4499 , w104 );
nor ( w4501 , w4500 , g1 );
nor ( w4502 , w4501 , g2 );
and ( w4503 , w4502 , g13 );
not ( w4504 , w4503 );
and ( w4505 , w4504 , w4455 );
and ( w4506 , w4505 , g3 );
and ( w4507 , w4506 , w8860 );
and ( w4508 , w4507 , g11 );
not ( w4509 , w4508 );
and ( w4510 , w4509 , w3767 );
and ( w4511 , w4510 , g12 );
not ( w4512 , w4511 );
and ( w4513 , w4512 , g3 );
and ( w4514 , w4513 , w408 );
not ( w4515 , w4514 );
and ( w4516 , w4515 , w4285 );
nor ( w4517 , w4516 , g16 );
not ( w4518 , w4471 );
and ( w4519 , w4518 , w4517 );
and ( w4520 , w4519 , w8860 );
and ( w4521 , w4520 , g11 );
and ( w4522 , w4521 , w7997 );
not ( w4523 , w4522 );
and ( w4524 , w4523 , w3767 );
and ( w4525 , w4524 , g12 );
not ( w4526 , w4525 );
and ( w4527 , w4526 , g3 );
not ( w4528 , w4527 );
and ( w4529 , w4528 , w4285 );
nor ( w4530 , w4529 , g9 );
and ( w4531 , w4530 , w8828 );
nor ( w4532 , w4440 , w4531 );
not ( w4533 , w4415 );
and ( w4534 , w4533 , w4532 );
nor ( w4535 , w4349 , w4534 );
and ( w4536 , w4535 , g3 );
not ( w4537 , w4536 );
and ( w4538 , w4537 , w4285 );
nor ( w4539 , w4538 , g6 );
not ( w4540 , w643 );
and ( w4541 , w4540 , g3 );
and ( w4542 , w4541 , w8765 );
and ( w4543 , w4542 , w7997 );
and ( w4544 , w4543 , w7783 );
nor ( w4545 , w4539 , w4544 );
not ( w4546 , w4545 );
and ( w4547 , w4546 , w1653 );
not ( w4548 , w4544 );
and ( w4549 , w4285 , w4548 );
and ( w4550 , w527 , w8819 );
not ( w4551 , w4550 );
and ( w4552 , w4551 , w4285 );
not ( w4553 , w4552 );
and ( w4554 , w4553 , g11 );
nor ( w4555 , w4554 , g12 );
and ( w4556 , w4555 , w4285 );
nor ( w4557 , w4556 , g16 );
not ( w4558 , w4557 );
and ( w4559 , w4549 , w4558 );
not ( w4560 , w4559 );
and ( w4561 , w4560 , g11 );
and ( w4562 , w4561 , w7997 );
not ( w4563 , w4562 );
and ( w4564 , w4563 , w3767 );
and ( w4565 , w4564 , w8728 );
and ( w4566 , w4565 , w4285 );
nor ( w4567 , w4566 , g16 );
nor ( w4568 , w4547 , w4567 );
nor ( w4569 , w4568 , g13 );
and ( w4570 , w518 , g6 );
and ( w4571 , w4570 , w299 );
and ( w4572 , w4571 , g3 );
and ( w4573 , w4572 , w7997 );
not ( w4574 , w4573 );
and ( w4575 , w4574 , w4285 );
not ( w4576 , w4575 );
and ( w4577 , w4576 , w4338 );
and ( w4578 , w4577 , g6 );
and ( w4579 , w4578 , w1489 );
and ( w4580 , w4579 , g13 );
and ( w4581 , w4580 , g11 );
not ( w4582 , w4581 );
and ( w4583 , w4582 , w3767 );
not ( w4584 , w4583 );
and ( w4585 , w4584 , g10 );
and ( w4586 , w4338 , g14 );
and ( w4587 , w4586 , g15 );
nor ( w4588 , w4587 , w4542 );
nor ( w4589 , w4588 , g13 );
not ( w4590 , w4589 );
and ( w4591 , w4590 , w4285 );
not ( w4592 , w4591 );
and ( w4593 , w4592 , g6 );
and ( w4594 , w7934 , w4538 );
nor ( w4595 , w4594 , g13 );
and ( w4596 , w4375 , w8792 );
not ( w4597 , w4359 );
and ( w4598 , w4596 , w4597 );
and ( w4599 , w4598 , g14 );
and ( w4600 , w4599 , g13 );
and ( w4601 , w4600 , w104 );
nor ( w4602 , w4601 , g12 );
nor ( w4603 , w4602 , w4534 );
and ( w4604 , w4603 , g3 );
not ( w4605 , w4604 );
and ( w4606 , w4605 , w4285 );
not ( w4607 , w4595 );
and ( w4608 , w4607 , w4606 );
not ( w4609 , w4608 );
and ( w4610 , w4609 , w4338 );
and ( w4611 , w4610 , w8845 );
and ( w4612 , w4611 , g11 );
and ( w4613 , w4612 , w7783 );
and ( w4614 , w4613 , g3 );
nor ( w4615 , w4614 , g12 );
nor ( w4616 , w4615 , w4534 );
and ( w4617 , w4616 , g3 );
not ( w4618 , w4617 );
and ( w4619 , w4618 , w4285 );
not ( w4620 , w4593 );
and ( w4621 , w4620 , w4619 );
not ( w4622 , w4621 );
and ( w4623 , w4622 , g11 );
not ( w4624 , w4623 );
and ( w4625 , w4624 , w4285 );
nor ( w4626 , w4625 , g10 );
and ( w4627 , w4626 , w7783 );
and ( w4628 , w4627 , g3 );
nor ( w4629 , w4628 , g12 );
nor ( w4630 , w4629 , w4534 );
and ( w4631 , w4630 , g3 );
not ( w4632 , w4631 );
and ( w4633 , w4632 , w4285 );
not ( w4634 , w4585 );
and ( w4635 , w4634 , w4633 );
nor ( w4636 , w4635 , g2 );
and ( w4637 , w4636 , g3 );
nor ( w4638 , w4637 , g12 );
nor ( w4639 , w4638 , w4534 );
and ( w4640 , w4639 , g3 );
not ( w4641 , w4640 );
and ( w4642 , w4641 , w4285 );
not ( w4643 , w4569 );
and ( w4644 , w4643 , w4642 );
not ( w4645 , w4644 );
and ( w4646 , w4645 , g11 );
and ( w4647 , w4646 , w7997 );
not ( w4648 , w4647 );
and ( w4649 , w4648 , w3767 );
not ( w4650 , w4649 );
and ( w4651 , w4650 , g10 );
not ( w4652 , w4651 );
and ( w4653 , w4652 , w4633 );
nor ( w4654 , w4653 , g2 );
and ( w4655 , w4654 , g3 );
nor ( w4656 , w4655 , g12 );
nor ( w4657 , w4656 , w4534 );
and ( w4658 , w4657 , g3 );
not ( w4659 , w4658 );
and ( w4660 , w4659 , w4285 );
not ( w4661 , w4342 );
and ( w4662 , w4661 , w4660 );
not ( w4663 , w4662 );
and ( w4664 , w4663 , w33 );
not ( w4665 , w4664 );
and ( w4666 , w4665 , w4633 );
nor ( w4667 , w4666 , g2 );
and ( w4668 , w4667 , g3 );
nor ( w4669 , w4668 , g12 );
nor ( w4670 , w4669 , w4534 );
and ( w4671 , w4670 , g3 );
not ( w4672 , w4671 );
and ( w4673 , w4672 , w4285 );
not ( w4674 , w4321 );
and ( w4675 , w4674 , w4673 );
and ( w4676 , w4675 , w8728 );
nor ( w4677 , w4676 , w4534 );
and ( w4678 , w4677 , w8792 );
and ( w4679 , w4678 , g3 );
not ( w4680 , w4679 );
and ( w4681 , w4680 , w4285 );
not ( w4682 , w3909 );
and ( w4683 , w4682 , w4681 );
not ( w4684 , w4683 );
and ( w4685 , w4684 , g6 );
nor ( w4686 , w4685 , w4302 );
not ( w4687 , w4686 );
and ( w4688 , w4687 , g11 );
not ( w4689 , w4688 );
and ( w4690 , w4689 , w4285 );
not ( w4691 , w4318 );
and ( w4692 , w4690 , w4691 );
not ( w4693 , w4692 );
and ( w4694 , w4693 , w4338 );
and ( w4695 , w4694 , g2 );
not ( w4696 , w4695 );
and ( w4697 , w4696 , w4673 );
and ( w4698 , w4697 , w8728 );
nor ( w4699 , w4698 , w4534 );
nor ( w4700 , w3702 , w4699 );
nor ( w4701 , w3698 , w4700 );
not ( w4702 , w4701 );
and ( w4703 , w4702 , w4285 );
and ( w4704 , w5332 , w4703 );
nor ( w4705 , w4704 , g6 );
and ( w4706 , w4705 , g11 );
and ( w4707 , w4706 , g14 );
and ( w4708 , w4707 , g15 );
and ( w4709 , w4708 , w4338 );
not ( w4710 , w4709 );
and ( w4711 , w4710 , g13 );
nor ( w4712 , w4711 , w4700 );
not ( w4713 , w4712 );
and ( w4714 , w4713 , w4285 );
not ( w4715 , w3676 );
and ( w4716 , w4715 , w4714 );
and ( w4717 , w4716 , g13 );
nor ( w4718 , w4717 , w4700 );
not ( w4719 , w4718 );
and ( w4720 , w3692 , w4719 );
nor ( w4721 , w4720 , g1 );
and ( w4722 , w4721 , g3 );
not ( w4723 , w4722 );
and ( w4724 , w4723 , g13 );
nor ( w4725 , w4724 , w4700 );
not ( w4726 , w4725 );
and ( w4727 , w4726 , w4285 );
and ( w4728 , w4572 , w8728 );
and ( w4729 , w4728 , w7997 );
and ( w4730 , w4729 , g13 );
not ( w4731 , w4730 );
and ( w4732 , w4731 , w4727 );
nor ( w4733 , w4732 , g1 );
and ( w4734 , w4733 , w8828 );
not ( w4735 , w4734 );
and ( w4736 , w4727 , w4735 );
not ( w4737 , w4736 );
and ( w4738 , w4737 , g6 );
and ( w4739 , w4738 , w7783 );
not ( w4740 , w4739 );
and ( w4741 , w4740 , w4727 );
not ( w4742 , w4741 );
and ( w4743 , w4742 , g11 );
not ( w4744 , w4743 );
and ( w4745 , w4744 , w4727 );
and ( w4746 , w8828 , w4745 );
nor ( w4747 , w4746 , g3 );
and ( w4748 , w4747 , w8860 );
and ( w4749 , w4748 , g10 );
and ( w4750 , w4749 , w8837 );
and ( w4751 , w4750 , g8 );
and ( w4752 , w4751 , w8845 );
and ( w4753 , w4752 , w4100 );
not ( w4754 , w4753 );
and ( w4755 , w4754 , w4745 );
not ( w4756 , w4755 );
and ( w4757 , w4756 , g14 );
and ( w4758 , w4757 , g15 );
not ( w4759 , w4758 );
and ( w4760 , w4759 , w4745 );
nor ( w4761 , w4760 , g9 );
and ( w4762 , w4761 , w7783 );
not ( w4763 , w4762 );
and ( w4764 , w4763 , w4745 );
nor ( w4765 , w4764 , g13 );
not ( w4766 , w4765 );
and ( w4767 , w4766 , w4745 );
not ( w4768 , w4746 );
and ( w4769 , w4768 , g6 );
not ( w4770 , w4769 );
and ( w4771 , w4770 , w4745 );
not ( w4772 , w4771 );
and ( w4773 , w4772 , g10 );
not ( w4774 , w4773 );
and ( w4775 , w4774 , w4745 );
nor ( w4776 , w4775 , g9 );
and ( w4777 , w4776 , g14 );
and ( w4778 , w4777 , g15 );
not ( w4779 , w4778 );
and ( w4780 , w4779 , w4745 );
not ( w4781 , w4780 );
and ( w4782 , w4781 , g11 );
not ( w4783 , w4782 );
and ( w4784 , w4783 , w4745 );
not ( w4785 , w4784 );
and ( w4786 , w4785 , g13 );
not ( w4787 , w4786 );
and ( w4788 , w4787 , w4745 );
not ( w4789 , w4788 );
and ( w4790 , w4789 , g2 );
not ( w4791 , w4790 );
and ( w4792 , w4791 , w4745 );
and ( t_8 , w4767 , w4792 );
nor ( w4793 , g1 , g10 );
nor ( w4794 , w4793 , g6 );
and ( w4795 , w4794 , g9 );
not ( w4796 , w4795 );
and ( w4797 , w4796 , g9 );
and ( w4798 , w2897 , g12 );
and ( w4799 , w4798 , w8382 );
and ( w4800 , w4799 , g14 );
and ( w4801 , w4800 , g3 );
and ( w4802 , w4801 , g9 );
and ( w4803 , w4802 , w8860 );
and ( w4804 , w4803 , w8837 );
and ( w4805 , w4804 , w8730 );
not ( w4806 , w4805 );
and ( w4807 , w4806 , g2 );
and ( w4808 , w1 , g9 );
and ( w4809 , w1845 , w8765 );
and ( w4810 , w4809 , w8742 );
and ( w4811 , w8769 , g6 );
and ( w4812 , w4810 , w4811 );
and ( w4813 , w4812 , w8792 );
nor ( w4814 , w4813 , g7 );
and ( w4815 , w4814 , w8860 );
and ( w4816 , w4815 , w8769 );
not ( w4817 , w4816 );
and ( w4818 , w4817 , g2 );
and ( w4819 , w1429 , w4818 );
and ( w4820 , w4819 , w8792 );
and ( w4821 , w4820 , g6 );
and ( w4822 , w4821 , g3 );
and ( w4823 , w4822 , g4 );
not ( w4824 , w2039 );
and ( w4825 , w408 , w4824 );
and ( w4826 , w4825 , w8860 );
and ( w4827 , w4826 , w526 );
nor ( w4828 , w44 , g4 );
and ( w4829 , w4828 , w8735 );
and ( w4830 , w4829 , w8765 );
nor ( w4831 , w4830 , g2 );
and ( w4832 , w4831 , w8845 );
and ( w4833 , w4832 , w8792 );
nor ( w4834 , w4449 , w4833 );
nor ( w4835 , w4834 , g1 );
and ( w4836 , w4835 , g9 );
nor ( w4837 , w4833 , g1 );
nor ( w4838 , w4837 , g2 );
and ( w4839 , w4838 , w8845 );
and ( w4840 , w4839 , w104 );
and ( w4841 , w4840 , w7783 );
not ( w4842 , w4837 );
and ( w4843 , w4842 , w4841 );
and ( w4844 , w4843 , w8845 );
and ( w4845 , w4844 , w7783 );
nor ( w4846 , g6 , w4845 );
not ( w4847 , w4846 );
and ( w4848 , w4847 , g1 );
and ( w4849 , g3 , g1 );
and ( w4850 , w1489 , w4849 );
not ( w4851 , w4850 );
and ( w4852 , w4851 , g3 );
not ( w4853 , w4852 );
and ( w4854 , w4853 , g1 );
and ( w4855 , w561 , w8769 );
and ( w4856 , w4855 , w8742 );
and ( w4857 , w3736 , w4880 );
and ( w4858 , w4857 , w408 );
nor ( w4859 , g9 , w4858 );
and ( w4860 , w4859 , g16 );
not ( w4861 , w4860 );
and ( w4862 , w4861 , g4 );
nor ( w4863 , w4862 , w381 );
nor ( w4864 , w4863 , g1 );
nor ( w4865 , w4864 , g11 );
nor ( w4866 , w4865 , g2 );
nor ( w4867 , w4854 , w4866 );
not ( w4868 , w4867 );
and ( w4869 , w4868 , g6 );
and ( w4870 , w6851 , w1751 );
and ( w4871 , w4870 , g9 );
and ( w4872 , w4871 , w104 );
and ( w4873 , w104 , w8765 );
nor ( w4874 , w4872 , w4873 );
not ( w4875 , w4874 );
and ( w4876 , w4875 , g1 );
nor ( w4877 , w297 , g3 );
not ( w4878 , w4877 );
and ( w4879 , w4878 , w408 );
not ( w4880 , w4856 );
and ( w4881 , w4879 , w4880 );
nor ( w4882 , w4881 , w381 );
not ( w4883 , w4882 );
and ( w4884 , w4883 , g4 );
nor ( w4885 , g9 , w4884 );
and ( w4886 , w1864 , w8769 );
and ( w4887 , w4886 , w8742 );
and ( w4888 , w4887 , w8845 );
and ( w4889 , w4888 , w8837 );
and ( w4890 , w4889 , g13 );
not ( w4891 , w4890 );
and ( w4892 , w4885 , w4891 );
nor ( w4893 , w4892 , g2 );
and ( w4894 , w4893 , w8845 );
not ( w4895 , w4894 );
and ( w4896 , w4895 , g16 );
not ( w4897 , w4896 );
and ( w4898 , w4897 , w4833 );
and ( w4899 , w4898 , g10 );
and ( w4900 , g2 , g9 );
and ( w4901 , w1651 , g6 );
not ( w4902 , w4901 );
and ( w4903 , w4902 , g6 );
not ( w4904 , w4903 );
and ( w4905 , w4900 , w4904 );
and ( w4906 , w4905 , g6 );
not ( w4907 , w4906 );
and ( w4908 , w4907 , g1 );
not ( w4909 , w4908 );
and ( w4910 , w4909 , w8882 );
and ( w4911 , w4910 , g6 );
and ( w4912 , g1 , g9 );
and ( w4913 , w4912 , w8845 );
and ( w4914 , w4913 , w400 );
nor ( w4915 , w4911 , w4914 );
not ( w4916 , w4915 );
and ( w4917 , w4916 , g3 );
nor ( w4918 , w4906 , w4914 );
nor ( w4919 , w4918 , g3 );
not ( w4920 , w4919 );
and ( w4921 , w4920 , g1 );
not ( w4922 , w4921 );
and ( w4923 , w4922 , w8882 );
nor ( w4924 , w4917 , w4923 );
not ( w4925 , w4924 );
and ( w4926 , w4925 , g9 );
not ( w4927 , w4926 );
and ( w4928 , w4927 , g9 );
not ( w4929 , w1521 );
and ( w4930 , w4929 , g9 );
nor ( w4931 , w4930 , g10 );
nor ( w4932 , w4931 , g10 );
and ( w4933 , w4932 , w8845 );
and ( w4934 , w4928 , w4933 );
nor ( w4935 , w4934 , w4873 );
not ( w4936 , w4935 );
and ( w4937 , w4936 , g1 );
and ( w4938 , w3679 , g4 );
not ( w4939 , w1395 );
and ( w4940 , w4939 , w361 );
and ( w4941 , w4940 , g5 );
and ( w4942 , w4941 , g7 );
and ( w4943 , w4942 , w8730 );
and ( w4944 , w4943 , g4 );
nor ( w4945 , w4944 , g3 );
and ( w4946 , w4945 , g5 );
and ( w4947 , w4946 , g7 );
and ( w4948 , w4947 , w8730 );
and ( w4949 , w4948 , g4 );
nor ( w4950 , w4949 , g6 );
nor ( w4951 , w4950 , g6 );
not ( w4952 , w4951 );
and ( w4953 , w4952 , w361 );
nor ( w4954 , w4953 , g9 );
nor ( w4955 , w4954 , g6 );
and ( w4956 , w4955 , g10 );
and ( w4957 , w4956 , g9 );
and ( w4958 , w4957 , w4849 );
not ( w4959 , w4958 );
and ( w4960 , w4959 , g3 );
not ( w4961 , w2190 );
and ( w4962 , w4960 , w4961 );
nor ( w4963 , w4962 , w1588 );
and ( w4964 , w4963 , w7783 );
and ( w4965 , w4964 , w8845 );
and ( w4966 , w8860 , w104 );
and ( w4967 , w4966 , w8792 );
and ( w4968 , w4967 , g10 );
not ( w4969 , w4934 );
and ( w4970 , w4969 , g9 );
not ( w4971 , w4970 );
and ( w4972 , w4971 , g1 );
and ( w4973 , w4972 , w8730 );
and ( w4974 , w4973 , w104 );
nor ( w4975 , w4974 , w4967 );
nor ( w4976 , w4975 , g4 );
and ( w4977 , w4976 , w8730 );
nor ( w4978 , w1489 , w4977 );
nor ( w4979 , w4978 , g4 );
and ( w4980 , w4979 , w8730 );
nor ( w4981 , w4968 , w4980 );
and ( w4982 , w8845 , w4981 );
nor ( w4983 , w4982 , g2 );
and ( w4984 , w4983 , w8792 );
and ( w4985 , w4984 , g10 );
nor ( w4986 , w4985 , w4980 );
nor ( w4987 , w4986 , g4 );
nor ( w4988 , w4965 , w4987 );
not ( w4989 , w4988 );
and ( w4990 , w4989 , g10 );
nor ( w4991 , w4990 , w4980 );
nor ( w4992 , w4991 , g4 );
nor ( w4993 , g6 , w4992 );
not ( w4994 , w4993 );
and ( w4995 , w4994 , g1 );
nor ( w4996 , w4995 , w4987 );
not ( w4997 , w4996 );
and ( w4998 , w4997 , g10 );
nor ( w4999 , w4998 , w4980 );
nor ( w5000 , w4999 , g4 );
and ( w5001 , w5000 , w7783 );
nor ( w5002 , w4938 , w5001 );
not ( w5003 , w4937 );
and ( w5004 , w5003 , w5002 );
not ( w5005 , w4899 );
and ( w5006 , w5005 , w5004 );
and ( w5007 , w5006 , w8837 );
nor ( w5008 , w5007 , g2 );
not ( w5009 , w5008 );
and ( w5010 , w5009 , g13 );
not ( w5011 , w4876 );
and ( w5012 , w5011 , w5010 );
not ( w5013 , w5012 );
and ( w5014 , w5013 , g10 );
not ( w5015 , w5014 );
and ( w5016 , w5015 , w5004 );
not ( w5017 , w5016 );
and ( w5018 , w5017 , w104 );
and ( w5019 , w5018 , w8845 );
and ( w5020 , w5019 , g4 );
nor ( w5021 , w5020 , w5001 );
not ( w5022 , w4869 );
and ( w5023 , w5022 , w5021 );
not ( w5024 , w5023 );
and ( w5025 , w5024 , g4 );
nor ( w5026 , w5025 , w5001 );
nor ( w5027 , w5026 , g2 );
not ( w5028 , w5027 );
and ( w5029 , w5028 , g13 );
and ( w5030 , w41 , w5033 );
nor ( w5031 , w4848 , w5030 );
nor ( w5032 , w5031 , g9 );
not ( w5033 , w5029 );
and ( w5034 , w5032 , w5033 );
and ( w5035 , w5034 , w7783 );
nor ( w5036 , w4836 , w5035 );
nor ( w5037 , w5036 , w5029 );
and ( w5038 , w5037 , w7783 );
nor ( w5039 , w2441 , w5038 );
not ( w5040 , w5039 );
and ( w5041 , w5040 , g6 );
nor ( w5042 , w5041 , w471 );
not ( w5043 , w5042 );
and ( w5044 , w5043 , w408 );
nor ( w5045 , w4827 , w5044 );
not ( w5046 , w4823 );
and ( w5047 , w5046 , w5045 );
not ( w5048 , w4808 );
and ( w5049 , w5048 , w5047 );
and ( w5050 , w5049 , w5151 );
not ( w5051 , w5050 );
and ( w5052 , w5051 , g4 );
and ( w5053 , w7070 , w1588 );
and ( w5054 , w5053 , g3 );
nor ( w5055 , w5054 , w27 );
nor ( w5056 , w5055 , g2 );
and ( w5057 , w5056 , w8860 );
nor ( w5058 , w5057 , g12 );
nor ( w5059 , w5058 , g2 );
and ( w5060 , w5059 , w8860 );
nor ( w5061 , w5060 , g13 );
and ( w5062 , w5061 , g11 );
and ( w5063 , w5062 , w7934 );
nor ( w5064 , w5063 , g1 );
nor ( w5065 , g2 , w5064 );
not ( w5066 , w5065 );
and ( w5067 , w5066 , g3 );
not ( w5068 , w5067 );
and ( w5069 , w5068 , g3 );
nor ( w5070 , w5069 , g6 );
nor ( w5071 , w5070 , g12 );
and ( w5072 , w5071 , w8819 );
nor ( w5073 , w5072 , g4 );
not ( w5074 , w5073 );
and ( w5075 , w5074 , g11 );
nor ( w5076 , w2075 , g3 );
and ( w5077 , w5076 , g4 );
and ( w5078 , w4570 , g7 );
and ( w5079 , w5078 , w270 );
not ( w5080 , w5079 );
and ( w5081 , w5080 , g7 );
nor ( w5082 , w5081 , g4 );
and ( w5083 , w5082 , g15 );
and ( w5084 , w5083 , w8730 );
nor ( w5085 , w5084 , w122 );
and ( w5086 , w5085 , w8730 );
not ( w5087 , w5086 );
and ( w5088 , w5087 , w291 );
and ( w5089 , w5088 , w2585 );
nor ( w5090 , w5089 , g3 );
and ( w5091 , w291 , g10 );
and ( w5092 , w5091 , w8769 );
and ( w5093 , w5092 , w8742 );
and ( w5094 , w5093 , g8 );
nor ( w5095 , w5094 , g5 );
and ( w5096 , w5095 , w8742 );
and ( w5097 , w5096 , g8 );
nor ( w5098 , w17 , g5 );
nor ( w5099 , w5097 , w5098 );
and ( w5100 , w5099 , w27 );
and ( w5101 , w5100 , w33 );
not ( w5102 , w5101 );
and ( w5103 , w5102 , w73 );
not ( w5104 , w5103 );
and ( w5105 , w5104 , g2 );
and ( w5106 , w5105 , w8765 );
nor ( w5107 , g4 , w5106 );
not ( w5108 , w5107 );
and ( w5109 , w5108 , g10 );
not ( w5110 , w5109 );
and ( w5111 , w5110 , w73 );
nor ( w5112 , w5111 , g3 );
and ( w5113 , w5112 , g2 );
not ( w5114 , w5113 );
and ( w5115 , w5114 , g2 );
and ( w5116 , w5115 , w8792 );
nor ( w5117 , w5116 , g9 );
nor ( w5118 , w5117 , g9 );
not ( w5119 , w5118 );
and ( w5120 , w5119 , g3 );
nor ( w5121 , w5120 , g1 );
not ( w5122 , w5090 );
and ( w5123 , w5122 , w5121 );
and ( w5124 , w5123 , w2585 );
nor ( w5125 , w5077 , w5124 );
and ( w5126 , w289 , w8742 );
and ( w5127 , w5126 , g5 );
and ( w5128 , w5127 , w8730 );
and ( w5129 , w5128 , g6 );
and ( w5130 , w5129 , w4184 );
and ( w5131 , w5130 , g4 );
nor ( w5132 , w5131 , g7 );
and ( w5133 , w5132 , g5 );
not ( w5134 , w5133 );
and ( w5135 , w5134 , w4418 );
not ( w5136 , w5135 );
and ( w5137 , w5136 , g4 );
not ( w5138 , w5137 );
and ( w5139 , w5138 , g6 );
not ( w5140 , w5125 );
and ( w5141 , w5140 , w5139 );
and ( w5142 , w5141 , w8735 );
nor ( w5143 , w5142 , g3 );
not ( w5144 , w5143 );
and ( w5145 , w5144 , w5121 );
and ( w5146 , w5145 , g2 );
and ( w5147 , w5146 , w2585 );
and ( w5148 , w5147 , w408 );
and ( w5149 , w5148 , w8730 );
nor ( w5150 , w5149 , g10 );
not ( w5151 , w5038 );
and ( w5152 , w5150 , w5151 );
not ( w5153 , w5152 );
and ( w5154 , w5153 , g6 );
and ( w5155 , w5154 , w8792 );
and ( w5156 , w5292 , w5155 );
nor ( w5157 , g9 , w471 );
nor ( w5158 , w1857 , g6 );
and ( w5159 , w5158 , w8792 );
and ( w5160 , w5159 , w8735 );
and ( w5161 , w5160 , w27 );
nor ( w5162 , g3 , w5161 );
not ( w5163 , w5162 );
and ( w5164 , w5163 , g2 );
and ( w5165 , w361 , w8728 );
and ( w5166 , w5165 , g7 );
and ( w5167 , w5166 , g11 );
not ( w5168 , w5167 );
and ( w5169 , w5164 , w5168 );
nor ( w5170 , w5169 , w122 );
and ( w5171 , w5170 , w8730 );
nor ( w5172 , w2711 , g7 );
nor ( w5173 , w5172 , g4 );
and ( w5174 , w5173 , w132 );
not ( w5175 , w5174 );
and ( w5176 , w5175 , g3 );
nor ( w5177 , w5176 , g9 );
nor ( w5178 , w5177 , g9 );
not ( w5179 , w5178 );
and ( w5180 , w5179 , g2 );
and ( w5181 , w5180 , w5336 );
and ( w5182 , w5181 , w8860 );
and ( w5183 , w5182 , w8765 );
and ( w5184 , w5183 , w8792 );
nor ( w5185 , w5184 , g9 );
nor ( w5186 , w5185 , g6 );
and ( w5187 , w5186 , g2 );
and ( w5188 , w5187 , w8860 );
and ( w5189 , w5188 , w8792 );
not ( w5190 , w5171 );
and ( w5191 , w5190 , w5189 );
nor ( w5192 , w5191 , g5 );
nor ( w5193 , w5192 , g4 );
and ( w5194 , w5193 , w241 );
nor ( w5195 , w5194 , g14 );
not ( w5196 , w5195 );
and ( w5197 , w5196 , w241 );
and ( w5198 , w5197 , w8860 );
nor ( w5199 , w5198 , g4 );
not ( w5200 , w5199 );
and ( w5201 , w5200 , w241 );
and ( w5202 , w5201 , w7997 );
nor ( w5203 , g6 , g14 );
and ( w5204 , w5203 , w8792 );
and ( w5205 , w5204 , w7783 );
nor ( w5206 , w5205 , w122 );
not ( w5207 , w5206 );
and ( w5208 , w5207 , w4833 );
nor ( w5209 , w5202 , w5208 );
nor ( w5210 , w5209 , g16 );
and ( w5211 , w5210 , g3 );
nor ( w5212 , w5161 , g4 );
nor ( w5213 , w5212 , g6 );
nor ( w5214 , w5211 , w5213 );
not ( w5215 , w5214 );
and ( w5216 , w5215 , g2 );
and ( w5217 , w5216 , w8860 );
nor ( w5218 , w5217 , g4 );
nor ( w5219 , w5218 , w5047 );
nor ( w5220 , w400 , w3679 );
not ( w5221 , w1515 );
and ( w5222 , w5220 , w5221 );
nor ( w5223 , w5222 , g1 );
and ( w5224 , w5219 , w5223 );
and ( w5225 , w5224 , g2 );
nor ( w5226 , w5225 , w5208 );
and ( w5227 , w5226 , w8828 );
nor ( w5228 , w5227 , g9 );
nor ( w5229 , w5228 , w381 );
nor ( w5230 , w5229 , g1 );
nor ( w5231 , w4900 , w5230 );
not ( w5232 , w5231 );
and ( w5233 , w5232 , g2 );
nor ( w5234 , w5233 , w5208 );
nor ( w5235 , w5234 , g6 );
nor ( w5236 , w5235 , w381 );
nor ( w5237 , w5236 , g1 );
not ( w5238 , w5157 );
and ( w5239 , w5238 , w5237 );
and ( w5240 , w5239 , w8845 );
and ( w5241 , w5240 , w8792 );
nor ( w5242 , w5156 , w5241 );
not ( w5243 , w4449 );
and ( w5244 , w5243 , w5242 );
nor ( w5245 , w5244 , g1 );
not ( w5246 , w5075 );
and ( w5247 , w5246 , w5245 );
nor ( w5248 , w5247 , w381 );
and ( w5249 , w8845 , w5248 );
and ( w5250 , w92 , g6 );
and ( w5251 , w5250 , g15 );
and ( w5252 , w5251 , g2 );
and ( w5253 , w5252 , w8742 );
nor ( w5254 , w5249 , w5253 );
nor ( w5255 , w5254 , g12 );
and ( w5256 , w8860 , g6 );
and ( w5257 , w5064 , w8845 );
and ( w5258 , w5257 , w7783 );
and ( w5259 , w5258 , w8860 );
nor ( w5260 , w5256 , w5259 );
nor ( w5261 , w5260 , g2 );
and ( w5262 , w5261 , w5245 );
nor ( w5263 , w290 , w5262 );
nor ( w5264 , w5263 , g9 );
nor ( w5265 , w5264 , g16 );
not ( w5266 , w4827 );
and ( w5267 , w5266 , g6 );
and ( w5268 , w5267 , g3 );
nor ( w5269 , w5268 , g2 );
nor ( w5270 , w5269 , g2 );
nor ( w5271 , w5270 , g4 );
and ( w5272 , w5271 , w8792 );
not ( w5273 , w5265 );
and ( w5274 , w5273 , w5272 );
and ( w5275 , w5274 , w8765 );
not ( w5276 , w5255 );
and ( w5277 , w5276 , w5275 );
nor ( w5278 , w5277 , g16 );
not ( w5279 , w5278 );
and ( w5280 , w5279 , w5272 );
nor ( w5281 , w5280 , g13 );
nor ( w5282 , w5281 , g9 );
and ( w5283 , w5282 , w5292 );
and ( w5284 , w5283 , w2687 );
not ( w5285 , w5284 );
and ( w5286 , w5285 , g11 );
not ( w5287 , w5286 );
and ( w5288 , w5287 , w5245 );
nor ( w5289 , w5288 , w381 );
not ( w5290 , w5289 );
and ( w5291 , w5290 , w5272 );
not ( w5292 , w5047 );
and ( w5293 , w5291 , w5292 );
nor ( w5294 , w1430 , w5293 );
nor ( w5295 , w5294 , g4 );
nor ( w5296 , w5052 , w5295 );
not ( w5297 , w5296 );
and ( w5298 , w5297 , w5245 );
not ( w5299 , w5298 );
and ( w5300 , w1588 , w5299 );
and ( w5301 , w4807 , w5685 );
nor ( w5302 , g1 , w5038 );
not ( w5303 , w5302 );
and ( w5304 , w5303 , g9 );
nor ( w5305 , w5304 , w5035 );
nor ( w5306 , w5305 , w5029 );
and ( w5307 , w5306 , w7783 );
nor ( w5308 , w5301 , w5307 );
and ( w5309 , w5308 , g13 );
nor ( w5310 , w4797 , w5309 );
and ( w5311 , w5310 , g1 );
nor ( w5312 , w4833 , w400 );
and ( w5313 , w6755 , w213 );
not ( w5314 , w5313 );
and ( w5315 , w5314 , g2 );
and ( w5316 , w5315 , w2585 );
and ( w5317 , w1473 , g2 );
and ( w5318 , w5317 , w8730 );
nor ( w5319 , w5318 , g8 );
nor ( w5320 , w5319 , g10 );
and ( w5321 , w7973 , g9 );
and ( w5322 , w5321 , g8 );
not ( w5323 , w5322 );
and ( w5324 , w5320 , w5323 );
nor ( w5325 , w5324 , w1347 );
nor ( w5326 , w5325 , g6 );
not ( w5327 , w5326 );
and ( w5328 , w5327 , g11 );
nor ( w5329 , w5328 , g6 );
and ( w5330 , w5329 , g2 );
nor ( w5331 , w5330 , w4833 );
not ( w5332 , w3695 );
and ( w5333 , w5332 , g2 );
nor ( w5334 , w5333 , g6 );
and ( w5335 , w5334 , w8792 );
not ( w5336 , w2847 );
and ( w5337 , w5336 , w5335 );
and ( w5338 , w5337 , w8845 );
and ( w5339 , w5338 , w8792 );
not ( w5340 , w5331 );
and ( w5341 , w5340 , w5339 );
and ( w5342 , w5341 , g13 );
nor ( w5343 , w5342 , g16 );
and ( w5344 , w5343 , w213 );
not ( w5345 , w5344 );
and ( w5346 , w5345 , w5237 );
not ( w5347 , w5346 );
and ( w5348 , w5347 , g13 );
not ( w5349 , w5316 );
and ( w5350 , w5349 , w5348 );
not ( w5351 , w5350 );
and ( w5352 , w5351 , g2 );
not ( w5353 , w2382 );
and ( w5354 , w5353 , g4 );
not ( w5355 , w5354 );
and ( w5356 , w5355 , w213 );
nor ( w5357 , w5356 , w5047 );
not ( w5358 , w5357 );
and ( w5359 , w5358 , g13 );
not ( w5360 , w5359 );
and ( w5361 , w5360 , g4 );
nor ( w5362 , w5361 , g16 );
nor ( w5363 , w5362 , g9 );
and ( w5364 , w5363 , w8792 );
and ( w5365 , g4 , w5364 );
and ( w5366 , w5365 , g6 );
and ( w5367 , w467 , w8792 );
nor ( w5368 , w5344 , w5047 );
not ( w5369 , w5368 );
and ( w5370 , w5369 , g13 );
not ( w5371 , w5370 );
and ( w5372 , w5367 , w5371 );
and ( w5373 , w5372 , w8765 );
nor ( w5374 , w5366 , w5373 );
and ( w5375 , w8742 , w27 );
and ( w5376 , w5375 , g8 );
and ( w5377 , w5376 , w17 );
nor ( w5378 , w5377 , g5 );
and ( w5379 , w5378 , w8735 );
and ( w5380 , w5379 , w8860 );
and ( w5381 , w5380 , w8742 );
nor ( w5382 , g1 , w5381 );
and ( w5383 , w5382 , w7783 );
and ( w5384 , w5383 , w13 );
nor ( w5385 , w5384 , g3 );
nor ( w5386 , w5385 , w5300 );
nor ( w5387 , g2 , w5386 );
nor ( w5388 , w5387 , g1 );
and ( w5389 , w5388 , w8765 );
and ( w5390 , w5389 , w8860 );
and ( w5391 , w5390 , w8735 );
and ( w5392 , w5391 , w8769 );
and ( w5393 , w5392 , w1244 );
and ( w5394 , w5393 , g10 );
nor ( w5395 , w5394 , g5 );
and ( w5396 , w5395 , w8735 );
and ( w5397 , w5396 , w8860 );
and ( w5398 , w5397 , g10 );
nor ( w5399 , w5398 , g7 );
nor ( w5400 , w5399 , g7 );
not ( w5401 , w5400 );
and ( w5402 , w5401 , g8 );
not ( w5403 , w5402 );
and ( w5404 , w5403 , g8 );
not ( w5405 , w5404 );
and ( w5406 , w5405 , g6 );
nor ( w5407 , w5092 , g5 );
and ( w5408 , w5407 , w8735 );
and ( w5409 , w5408 , g10 );
nor ( w5410 , w5409 , g7 );
nor ( w5411 , w5410 , g7 );
not ( w5412 , w765 );
and ( w5413 , w5412 , w27 );
nor ( w5414 , w5413 , g3 );
not ( w5415 , w5414 );
and ( w5416 , w5415 , g8 );
nor ( w5417 , g8 , w5300 );
nor ( w5418 , w5416 , w5417 );
nor ( w5419 , w5418 , w5300 );
and ( w5420 , w5419 , w8792 );
not ( w5421 , w5411 );
and ( w5422 , w5421 , w5420 );
and ( w5423 , w5422 , g8 );
nor ( w5424 , w5423 , w5417 );
not ( w5425 , w5424 );
and ( w5426 , w5425 , g2 );
nor ( w5427 , w1517 , w5307 );
nor ( w5428 , w5427 , w5300 );
and ( w5429 , w5428 , g6 );
not ( w5430 , w3679 );
and ( w5431 , w5430 , w213 );
not ( w5432 , w5431 );
and ( w5433 , w5432 , w5307 );
not ( w5434 , w5433 );
and ( w5435 , w5434 , g16 );
not ( w5436 , w5342 );
and ( w5437 , w5436 , w213 );
nor ( w5438 , w5437 , g6 );
and ( w5439 , w5438 , w5237 );
nor ( w5440 , w5439 , g16 );
nor ( w5441 , w5440 , g6 );
not ( w5442 , w5441 );
and ( w5443 , w5442 , g13 );
and ( w5444 , w5443 , w8837 );
nor ( w5445 , w5444 , g1 );
not ( w5446 , w5435 );
and ( w5447 , w5446 , w5445 );
and ( w5448 , w5447 , w8845 );
not ( w5449 , w5448 );
and ( w5450 , w5449 , g13 );
and ( w5451 , w5450 , w8837 );
nor ( w5452 , w5451 , g1 );
nor ( w5453 , w241 , w5452 );
nor ( w5454 , w5453 , g6 );
nor ( w5455 , w5429 , w5454 );
nor ( w5456 , w5455 , g1 );
and ( w5457 , w5426 , w5456 );
nor ( w5458 , g4 , w5457 );
not ( w5459 , w5458 );
and ( w5460 , w5459 , w400 );
not ( w5461 , w3192 );
and ( w5462 , w5461 , w27 );
and ( w5463 , w5462 , g8 );
and ( w5464 , w5463 , w17 );
nor ( w5465 , w5464 , g3 );
and ( w5466 , w5465 , g8 );
and ( w5467 , w5466 , w8769 );
and ( w5468 , w5467 , w8742 );
and ( w5469 , w5468 , w8860 );
nor ( w5470 , w5469 , g2 );
and ( w5471 , w5470 , w5685 );
nor ( w5472 , w5460 , w5471 );
nor ( w5473 , w5472 , g6 );
and ( w5474 , w5473 , w5456 );
nor ( w5475 , w5406 , w5474 );
nor ( w5476 , w5475 , g9 );
and ( w5477 , w5476 , w5685 );
and ( w5478 , w5477 , w5456 );
and ( w5479 , w5478 , g6 );
nor ( w5480 , g9 , w5370 );
and ( w5481 , w5480 , w8845 );
and ( w5482 , w5481 , w5685 );
and ( w5483 , w5482 , g4 );
and ( w5484 , g10 , g13 );
and ( w5485 , w5484 , w213 );
and ( w5486 , w5256 , g3 );
and ( w5487 , w5739 , w361 );
and ( w5488 , w5487 , w8860 );
nor ( w5489 , w5486 , w5488 );
nor ( w5490 , w5489 , w5253 );
nor ( w5491 , w5490 , g12 );
not ( w5492 , w5491 );
and ( w5493 , w5492 , g2 );
nor ( w5494 , w5493 , g13 );
nor ( w5495 , w5494 , w5047 );
nor ( w5496 , w5495 , w381 );
not ( w5497 , w5496 );
and ( w5498 , w5497 , g2 );
and ( w5499 , w5498 , g6 );
and ( w5500 , w5 , g10 );
nor ( w5501 , w5500 , g5 );
and ( w5502 , w5501 , w8735 );
and ( w5503 , w5502 , g10 );
nor ( w5504 , w5503 , g7 );
and ( w5505 , w5504 , g8 );
nor ( w5506 , w5505 , g7 );
and ( w5507 , w5506 , g8 );
not ( w5508 , w5507 );
and ( w5509 , w5508 , w472 );
and ( w5510 , w5167 , w8730 );
and ( w5511 , w5510 , g15 );
and ( w5512 , w5511 , w8769 );
and ( w5513 , w5512 , w7934 );
not ( w5514 , w5513 );
and ( w5515 , w5509 , w5514 );
nor ( w5516 , w5515 , g13 );
nor ( w5517 , w5516 , w5370 );
and ( w5518 , w5517 , w8845 );
and ( w5519 , w5518 , g2 );
and ( w5520 , w5519 , w8860 );
nor ( w5521 , w5520 , g16 );
nor ( w5522 , w5521 , g9 );
and ( w5523 , w5522 , w8792 );
nor ( w5524 , w5499 , w5523 );
not ( w5525 , w5524 );
and ( w5526 , w5525 , g2 );
and ( w5527 , w5526 , w8860 );
nor ( w5528 , w5527 , g16 );
nor ( w5529 , w5528 , g9 );
not ( w5530 , w5529 );
and ( w5531 , w5530 , g11 );
nor ( w5532 , w5531 , g1 );
not ( w5533 , w5485 );
and ( w5534 , w5533 , w5532 );
and ( w5535 , w5534 , g6 );
nor ( w5536 , w5535 , w5523 );
and ( w5537 , w1984 , w8860 );
not ( w5538 , w5537 );
and ( w5539 , w5538 , w17 );
nor ( w5540 , w5539 , g3 );
and ( w5541 , w5540 , w8769 );
nor ( w5542 , w5541 , g8 );
nor ( w5543 , w5542 , g8 );
not ( w5544 , w5543 );
and ( w5545 , w5544 , g2 );
not ( w5546 , w15 );
and ( w5547 , w5546 , w17 );
nor ( w5548 , w5547 , g8 );
and ( w5549 , w5548 , w8769 );
not ( w5550 , w5549 );
and ( w5551 , w5545 , w5550 );
and ( w5552 , w8710 , w5551 );
and ( w5553 , w5552 , w5685 );
nor ( w5554 , w5553 , w2022 );
and ( w5555 , w3190 , w59 );
and ( w5556 , w5555 , w17 );
nor ( w5557 , w5556 , g5 );
and ( w5558 , w5557 , g10 );
not ( w5559 , w5558 );
and ( w5560 , w5559 , w27 );
nor ( w5561 , w5560 , g3 );
not ( w5562 , w5561 );
and ( w5563 , w5562 , g8 );
not ( w5564 , w5563 );
and ( w5565 , w5564 , g8 );
and ( w5566 , w5565 , w8742 );
not ( w5567 , w5566 );
and ( w5568 , w5567 , g2 );
and ( w5569 , w5568 , w8792 );
not ( w5570 , w5569 );
and ( w5571 , w5570 , g2 );
nor ( w5572 , w5571 , g9 );
and ( w5573 , w5572 , w8792 );
not ( w5574 , w5554 );
and ( w5575 , w5574 , w5573 );
and ( w5576 , w5575 , g6 );
nor ( w5577 , w5576 , w472 );
nor ( w5578 , w290 , w519 );
and ( w5579 , w1 , w8860 );
not ( w5580 , w5579 );
and ( w5581 , w5580 , g2 );
nor ( w5582 , w5578 , w5581 );
and ( w5583 , w5582 , w8792 );
not ( w5584 , w5577 );
and ( w5585 , w5584 , w5583 );
nor ( w5586 , w5479 , w5474 );
and ( w5587 , w8765 , w5586 );
not ( w5588 , w5587 );
and ( w5589 , w5588 , w5456 );
and ( w5590 , w5585 , w5589 );
not ( w5591 , w5536 );
and ( w5592 , w5591 , w5590 );
and ( w5593 , w5592 , g2 );
nor ( w5594 , w3287 , g2 );
and ( w5595 , w5594 , w5589 );
and ( w5596 , w5595 , w4833 );
nor ( w5597 , w5596 , g6 );
not ( w5598 , w5597 );
and ( w5599 , w5598 , g10 );
not ( w5600 , w5599 );
and ( w5601 , w5600 , g10 );
nor ( w5602 , w5601 , g7 );
nor ( w5603 , w5602 , g7 );
nor ( w5604 , w5603 , g2 );
and ( w5605 , w5604 , w8860 );
and ( w5606 , w5605 , w8765 );
and ( w5607 , w5606 , w5589 );
nor ( w5608 , w5593 , w5607 );
and ( w5609 , w5608 , w8828 );
nor ( w5610 , w5609 , g9 );
not ( w5611 , w5610 );
and ( w5612 , w5611 , g11 );
not ( w5613 , w5612 );
and ( w5614 , w5613 , w5589 );
nor ( w5615 , w5483 , w5614 );
nor ( w5616 , w5615 , g9 );
and ( w5617 , w5616 , w5589 );
nor ( w5618 , w5479 , w5617 );
not ( w5619 , w5618 );
and ( w5620 , w5619 , g4 );
nor ( w5621 , w5620 , w5614 );
nor ( w5622 , w5621 , g9 );
not ( w5623 , w5374 );
and ( w5624 , w5623 , w5622 );
nor ( w5625 , w5624 , w5614 );
nor ( w5626 , w5625 , g9 );
nor ( w5627 , w2086 , w5626 );
not ( w5628 , w5627 );
and ( w5629 , w5628 , w5589 );
nor ( w5630 , w5352 , w5629 );
and ( w5631 , w5630 , g13 );
and ( w5632 , w5631 , w8828 );
not ( w5633 , w1517 );
and ( w5634 , w5633 , w5343 );
not ( w5635 , w5634 );
and ( w5636 , w5635 , g2 );
nor ( w5637 , w5636 , w5629 );
and ( w5638 , w5637 , g13 );
and ( w5639 , w5638 , w213 );
nor ( w5640 , w5639 , g1 );
and ( w5641 , w5640 , w5685 );
and ( w5642 , w5641 , g9 );
nor ( w5643 , w5642 , w5626 );
nor ( w5644 , w5632 , w5643 );
not ( w5645 , w5644 );
and ( w5646 , w5645 , g11 );
not ( w5647 , w5646 );
and ( w5648 , w5647 , w5589 );
not ( w5649 , w5312 );
and ( w5650 , w5649 , w5648 );
nor ( w5651 , w5311 , w5650 );
nor ( w5652 , w5651 , g6 );
not ( w5653 , w5652 );
and ( w5654 , w5653 , g16 );
and ( w5655 , w2847 , g1 );
not ( w5656 , w5655 );
and ( w5657 , w5656 , g1 );
nor ( w5658 , w5657 , w5650 );
nor ( w5659 , w5654 , w5658 );
nor ( w5660 , w2022 , w5659 );
not ( w5661 , w5660 );
and ( w5662 , w5661 , w5648 );
nor ( w5663 , g6 , w5659 );
and ( w5664 , w5711 , g1 );
nor ( w5665 , w5662 , w5664 );
nor ( w5666 , w5665 , g2 );
and ( w5667 , w2382 , g6 );
and ( w5668 , w5667 , w4849 );
and ( w5669 , w5668 , g9 );
not ( w5670 , w5669 );
and ( w5671 , w5670 , g10 );
and ( w5672 , w5671 , g3 );
not ( w5673 , w5672 );
and ( w5674 , w5673 , g6 );
and ( w5675 , w5674 , g2 );
and ( w5676 , w5675 , g1 );
nor ( w5677 , w5676 , w5659 );
not ( w5678 , w5677 );
and ( w5679 , w5678 , g9 );
and ( w5680 , w5679 , g1 );
and ( w5681 , w5680 , g2 );
not ( w5682 , w5681 );
and ( w5683 , w5682 , g9 );
nor ( w5684 , w5683 , w5663 );
not ( w5685 , w5300 );
and ( w5686 , w5684 , w5685 );
and ( w5687 , w5686 , g2 );
and ( w5688 , w5687 , g6 );
nor ( w5689 , w5688 , w5659 );
and ( w5690 , w5664 , g9 );
and ( w5691 , g2 , w5711 );
and ( w5692 , w5691 , w8765 );
nor ( w5693 , w5690 , w5692 );
not ( w5694 , w5659 );
and ( w5695 , w5694 , g7 );
and ( w5696 , w5695 , w8769 );
nor ( w5697 , w5659 , g7 );
and ( w5698 , w5697 , g5 );
nor ( w5699 , w5696 , w5698 );
not ( w5700 , w5699 );
and ( w5701 , w5700 , g17 );
and ( w5702 , w5701 , g12 );
and ( w5703 , w5702 , w8382 );
and ( w5704 , w5703 , g14 );
and ( w5705 , w5704 , g3 );
and ( w5706 , w5705 , g9 );
and ( w5707 , w5706 , w8860 );
and ( w5708 , w5707 , g10 );
not ( w5709 , w5708 );
and ( w5710 , w5709 , g2 );
not ( w5711 , w5663 );
and ( w5712 , w5710 , w5711 );
nor ( w5713 , w5712 , w5659 );
and ( w5714 , w5713 , w8837 );
nor ( w5715 , w5714 , w5663 );
and ( w5716 , w5715 , g2 );
nor ( w5717 , w5716 , w5659 );
nor ( w5718 , w5693 , w5717 );
and ( w5719 , w5718 , g2 );
and ( w5720 , w5719 , g6 );
nor ( w5721 , w5720 , w5659 );
and ( w5722 , w5721 , w8828 );
nor ( w5723 , w5722 , w5663 );
and ( w5724 , w5723 , g1 );
and ( w5725 , w5724 , g2 );
not ( w5726 , w5725 );
and ( w5727 , w5726 , g13 );
nor ( w5728 , w5727 , w5663 );
not ( w5729 , w5689 );
and ( w5730 , w5729 , w5728 );
and ( w5731 , w5730 , g1 );
nor ( w5732 , w5731 , w5648 );
not ( w5733 , w5732 );
and ( w5734 , w5733 , g2 );
nor ( t_9 , w5666 , w5734 );
nor ( w5735 , w468 , g6 );
not ( w5736 , w5735 );
and ( w5737 , w5736 , g4 );
and ( w5738 , w1845 , g3 );
not ( w5739 , w663 );
and ( w5740 , w5739 , g6 );
and ( w5741 , w5740 , w361 );
and ( w5742 , w5741 , w8792 );
nor ( w5743 , w5738 , w5742 );
not ( w5744 , w5743 );
and ( w5745 , w5744 , g2 );
and ( w5746 , w5745 , g6 );
and ( w5747 , w467 , w8735 );
not ( w5748 , w5747 );
and ( w5749 , w5748 , g4 );
and ( w5750 , w660 , w8730 );
nor ( w5751 , w5750 , w122 );
not ( w5752 , w5751 );
and ( w5753 , w5752 , w1613 );
nor ( w5754 , w5753 , g10 );
and ( w5755 , w5754 , g7 );
and ( w5756 , w5755 , w8769 );
and ( w5757 , w92 , g5 );
nor ( w5758 , w5757 , w1613 );
and ( w5759 , w92 , w8742 );
not ( w5760 , w5759 );
and ( w5761 , w5758 , w5760 );
nor ( w5762 , w5761 , g6 );
nor ( w5763 , w5762 , g6 );
nor ( w5764 , w5763 , g4 );
nor ( w5765 , w5764 , g4 );
nor ( w5766 , w5765 , g3 );
nor ( w5767 , w5766 , g10 );
and ( w5768 , w6688 , g5 );
nor ( w5769 , w5768 , w1613 );
nor ( w5770 , w123 , g15 );
and ( w5771 , g7 , w8730 );
not ( w5772 , w5770 );
and ( w5773 , w5772 , w5771 );
nor ( w5774 , w5773 , g10 );
nor ( w5775 , w5774 , w216 );
and ( w5776 , w5775 , w8792 );
and ( w5777 , w5776 , w8860 );
and ( w5778 , w5777 , w8735 );
not ( w5779 , w5769 );
and ( w5780 , w5779 , w5778 );
not ( w5781 , w5780 );
and ( w5782 , w5781 , g7 );
nor ( w5783 , w5782 , g4 );
and ( w5784 , w5783 , w361 );
nor ( w5785 , w5784 , g9 );
nor ( w5786 , w5785 , g1 );
not ( w5787 , w5756 );
and ( w5788 , w5787 , w5786 );
nor ( w5789 , w5788 , g4 );
not ( w5790 , w5789 );
and ( w5791 , w5790 , w770 );
and ( w5792 , w5791 , w361 );
and ( w5793 , w5792 , w408 );
nor ( w5794 , w5793 , g9 );
nor ( w5795 , w5794 , g1 );
not ( w5796 , w5749 );
and ( w5797 , w5796 , w5795 );
and ( w5798 , w5797 , w690 );
and ( w5799 , w5798 , w8845 );
and ( w5800 , w5799 , w8765 );
and ( w5801 , g10 , w8168 );
and ( w5802 , w5801 , g14 );
and ( w5803 , w4833 , w5456 );
and ( w5804 , w5803 , w8860 );
nor ( w5805 , w1852 , w5804 );
nor ( w5806 , w5805 , g1 );
and ( w5807 , w5806 , w7783 );
nor ( w5808 , w5807 , g12 );
nor ( w5809 , w5808 , g6 );
and ( w5810 , w5809 , w8792 );
and ( w5811 , w6160 , w5810 );
not ( w5812 , w5811 );
and ( w5813 , w5812 , g13 );
nor ( w5814 , w5813 , g2 );
nor ( w5815 , w5814 , g11 );
and ( w5816 , w5815 , w8728 );
nor ( w5817 , w5816 , g6 );
and ( w5818 , w5817 , w8792 );
nor ( w5819 , g9 , g2 );
and ( w5820 , w5818 , w5819 );
nor ( w5821 , w5820 , g11 );
and ( w5822 , w5821 , w8728 );
nor ( w5823 , w5822 , g6 );
and ( w5824 , w5823 , w8765 );
and ( w5825 , w5824 , w8792 );
nor ( w5826 , w5800 , w5825 );
and ( w5827 , w5826 , w8837 );
and ( w5828 , w5827 , g16 );
nor ( w5829 , g14 , g10 );
and ( w5830 , w5829 , g15 );
and ( w5831 , w5830 , w8860 );
and ( w5832 , w5831 , g7 );
and ( w5833 , w5832 , w8769 );
and ( w5834 , w5833 , g2 );
not ( w5835 , w5834 );
and ( w5836 , w5835 , w471 );
not ( w5837 , w5836 );
and ( w5838 , w5837 , g11 );
nor ( w5839 , g10 , w1366 );
not ( w5840 , w5839 );
and ( w5841 , w5840 , w2669 );
and ( w5842 , w5841 , w8730 );
not ( w5843 , w5842 );
and ( w5844 , w5843 , w1588 );
and ( w5845 , w3471 , g9 );
and ( w5846 , w5845 , g17 );
and ( w5847 , w5846 , g15 );
and ( w5848 , w5847 , g14 );
and ( w5849 , w5848 , g16 );
not ( w5850 , w5849 );
and ( w5851 , w5850 , g11 );
and ( w5852 , w1544 , w8845 );
and ( w5853 , w5852 , w8730 );
and ( w5854 , w5853 , g17 );
and ( w5855 , w5854 , w8769 );
and ( w5856 , w5855 , w8765 );
and ( w5857 , w5856 , w8742 );
and ( w5858 , w5857 , w8860 );
and ( w5859 , w5858 , g2 );
and ( w5860 , w5859 , g12 );
and ( w5861 , w5860 , g15 );
and ( w5862 , w5861 , g14 );
and ( w5863 , w5862 , g16 );
nor ( w5864 , w5863 , g11 );
not ( w5865 , w5864 );
and ( w5866 , w5865 , w400 );
and ( w5867 , w5866 , w8735 );
and ( w5868 , w5867 , w8792 );
not ( w5869 , w5851 );
and ( w5870 , w5869 , w5868 );
not ( w5871 , w5870 );
and ( w5872 , w5871 , g13 );
not ( w5873 , w5872 );
and ( w5874 , w5873 , w400 );
and ( w5875 , w5874 , w8735 );
and ( w5876 , w5875 , w8792 );
nor ( w5877 , w5844 , w5876 );
not ( w5878 , w5877 );
and ( w5879 , w5878 , g2 );
nor ( w5880 , w5431 , g1 );
and ( w5881 , w5880 , w40 );
nor ( w5882 , w5881 , g16 );
nor ( w5883 , w5882 , g2 );
and ( w5884 , w5883 , w4833 );
not ( w5885 , w5884 );
and ( w5886 , w5885 , g11 );
nor ( w5887 , w5886 , g6 );
not ( w5888 , w5887 );
and ( w5889 , w5888 , g13 );
nor ( w5890 , w5889 , g1 );
and ( w5891 , w5890 , w104 );
nor ( w5892 , w5879 , w5891 );
nor ( w5893 , w5892 , g3 );
nor ( w5894 , w5893 , g16 );
and ( w5895 , w5894 , w213 );
nor ( w5896 , w5895 , g6 );
not ( w5897 , w5896 );
and ( w5898 , w5897 , g11 );
and ( w5899 , w5898 , g13 );
nor ( w5900 , w5899 , g6 );
and ( w5901 , w5900 , w8735 );
and ( w5902 , w5901 , w8792 );
and ( w5903 , w5902 , w8765 );
not ( w5904 , w5903 );
and ( w5905 , w5904 , w213 );
not ( w5906 , w2126 );
and ( w5907 , w5906 , g8 );
not ( w5908 , w5907 );
and ( w5909 , w5908 , w33 );
nor ( w5910 , w5909 , g7 );
and ( w5911 , w5910 , g10 );
not ( w5912 , w5911 );
and ( w5913 , w5912 , w17 );
nor ( w5914 , w5913 , g5 );
not ( w5915 , w5914 );
and ( w5916 , w5915 , g2 );
not ( w5917 , w5916 );
and ( w5918 , w5917 , g2 );
nor ( w5919 , w1260 , g2 );
not ( w5920 , w270 );
and ( w5921 , w5920 , g7 );
not ( w5922 , w5921 );
and ( w5923 , w5922 , w17 );
nor ( w5924 , w5923 , w1786 );
not ( w5925 , w5924 );
and ( w5926 , w5925 , g8 );
nor ( w5927 , w5926 , w489 );
nor ( w5928 , w5919 , w5927 );
and ( w5929 , w27 , w8765 );
and ( w5930 , w5929 , w8792 );
and ( w5931 , w5930 , w8769 );
nor ( w5932 , w5931 , g5 );
not ( w5933 , w5932 );
and ( w5934 , w5933 , g2 );
and ( w5935 , w5934 , w8742 );
not ( w5936 , w5935 );
and ( w5937 , w5936 , g2 );
and ( w5938 , w5937 , w8742 );
not ( w5939 , w5938 );
and ( w5940 , w5939 , g8 );
not ( w5941 , w5940 );
and ( w5942 , w5941 , g8 );
not ( w5943 , w5942 );
and ( w5944 , w5928 , w5943 );
and ( w5945 , w5944 , g10 );
and ( w5946 , w5945 , w33 );
nor ( w5947 , w5946 , w92 );
nor ( w5948 , w5947 , g4 );
and ( w5949 , w5948 , w8792 );
not ( w5950 , w5918 );
and ( w5951 , w5950 , w5949 );
and ( w5952 , w5951 , w381 );
not ( w5953 , w5952 );
and ( w5954 , w5953 , w213 );
nor ( w5955 , w5954 , g6 );
and ( w5956 , w5955 , w8735 );
nor ( w5957 , w5956 , g9 );
nor ( w5958 , w5957 , g1 );
nor ( w5959 , w5958 , g1 );
nor ( w5960 , w5959 , g4 );
and ( w5961 , w5960 , w8735 );
and ( w5962 , w5961 , w8845 );
nor ( w5963 , w5962 , g3 );
nor ( w5964 , w5963 , g1 );
nor ( w5965 , w5964 , g1 );
and ( w5966 , w5965 , w8845 );
and ( w5967 , w518 , w27 );
and ( w5968 , w5967 , w408 );
nor ( w5969 , w5966 , w5968 );
not ( w5970 , w5969 );
and ( w5971 , w5970 , w400 );
nor ( w5972 , w5322 , w1367 );
and ( w5973 , w5972 , w8730 );
and ( w5974 , w5973 , w8845 );
nor ( w5975 , w5974 , g10 );
not ( w5976 , w5975 );
and ( w5977 , w5976 , g14 );
and ( w5978 , w5977 , g15 );
and ( w5979 , w3679 , g8 );
and ( w5980 , w5979 , g9 );
and ( w5981 , w5980 , w8382 );
and ( w5982 , w3679 , w8767 );
and ( w5983 , w5982 , g17 );
nor ( w5984 , w5981 , w5983 );
and ( w5985 , w5984 , w213 );
nor ( w5986 , w5985 , g1 );
and ( w5987 , w5986 , w40 );
and ( w5988 , w5987 , w8735 );
and ( w5989 , w5988 , w8845 );
not ( w5990 , w5989 );
and ( w5991 , w5990 , g13 );
nor ( w5992 , w5991 , g2 );
and ( w5993 , w5992 , w8845 );
and ( w5994 , w5993 , w8735 );
and ( w5995 , w5994 , w8792 );
nor ( w5996 , w5978 , w5995 );
and ( w5997 , w5996 , w8828 );
not ( w5998 , w5997 );
and ( w5999 , w5998 , w4833 );
not ( w6000 , w5999 );
and ( w6001 , w6000 , g11 );
and ( w6002 , w6001 , g13 );
nor ( w6003 , w6002 , g6 );
and ( w6004 , w6003 , w7783 );
and ( w6005 , w6160 , w6004 );
nor ( w6006 , w5995 , g16 );
nor ( w6007 , w6006 , g6 );
and ( w6008 , w6007 , w7783 );
and ( w6009 , w6008 , w8735 );
nor ( w6010 , w6005 , w6009 );
and ( w6011 , w6010 , w8828 );
nor ( w6012 , w6011 , g2 );
and ( w6013 , w6012 , w4833 );
not ( w6014 , w6013 );
and ( w6015 , w6014 , g11 );
nor ( w6016 , w6015 , g3 );
not ( w6017 , w6016 );
and ( w6018 , w6017 , g13 );
nor ( w6019 , w6018 , g1 );
and ( w6020 , w6019 , w104 );
and ( w6021 , w6020 , w8735 );
not ( w6022 , w6021 );
and ( w6023 , w6022 , g13 );
and ( w6024 , w6023 , w8828 );
nor ( w6025 , w6024 , g6 );
and ( w6026 , w6025 , w8792 );
nor ( w6027 , w5971 , w6026 );
and ( w6028 , w6027 , g11 );
and ( w6029 , w2224 , g2 );
and ( w6030 , w1260 , w8845 );
nor ( w6031 , w6029 , w6030 );
nor ( w6032 , w6031 , g3 );
and ( w6033 , w6032 , w8765 );
not ( w6034 , w6028 );
and ( w6035 , w6034 , w6033 );
not ( w6036 , w6035 );
and ( w6037 , w6036 , g13 );
nor ( w6038 , w6037 , g6 );
nor ( w6039 , w6038 , g16 );
nor ( w6040 , w6039 , g3 );
nor ( w6041 , w6040 , g12 );
and ( w6042 , w92 , w8860 );
nor ( w6043 , w6042 , g1 );
and ( w6044 , w400 , g4 );
and ( w6045 , w6043 , w6044 );
nor ( w6046 , w6045 , w3736 );
nor ( w6047 , w5800 , g9 );
nor ( w6048 , w6047 , g1 );
and ( w6049 , w6048 , g2 );
and ( w6050 , w6049 , w8845 );
not ( w6051 , w6050 );
and ( w6052 , w6051 , g2 );
nor ( w6053 , w6052 , g3 );
and ( w6054 , w6053 , g5 );
and ( w6055 , w2687 , w8765 );
nor ( w6056 , w6055 , g9 );
nor ( w6057 , w6056 , g4 );
and ( w6058 , w6057 , w8845 );
and ( w6059 , w6058 , w59 );
nor ( w6060 , w6059 , g7 );
and ( w6061 , w512 , w7783 );
and ( w6062 , w6061 , w8845 );
and ( w6063 , w6062 , g7 );
nor ( w6064 , w213 , g1 );
and ( w6065 , w6064 , w8845 );
not ( w6066 , w6065 );
and ( w6067 , w6066 , g16 );
not ( w6068 , w6067 );
and ( w6069 , w6068 , w6009 );
and ( w6070 , g13 , w6069 );
and ( w6071 , w6070 , g11 );
and ( w6072 , w6071 , g7 );
and ( w6073 , w566 , g14 );
and ( w6074 , w6073 , g15 );
nor ( w6075 , w6074 , g13 );
not ( w6076 , w6075 );
and ( w6077 , w6076 , w5995 );
and ( w6078 , w6077 , w8769 );
and ( w6079 , w6078 , w59 );
and ( w6080 , w6079 , g12 );
and ( w6081 , w6080 , w1844 );
and ( w6082 , w6081 , w8828 );
nor ( w6083 , w6082 , g13 );
and ( w6084 , w519 , w8767 );
and ( w6085 , w6084 , w8845 );
and ( w6086 , w6085 , w59 );
and ( w6087 , w6086 , g10 );
and ( w6088 , w6087 , w8735 );
and ( w6089 , w6088 , g12 );
not ( w6090 , w6089 );
and ( w6091 , w6090 , w213 );
nor ( w6092 , w6091 , g6 );
and ( w6093 , w6092 , w7783 );
not ( w6094 , w6093 );
and ( w6095 , w6094 , g16 );
not ( w6096 , w6095 );
and ( w6097 , w6096 , w6009 );
and ( w6098 , w6097 , w8792 );
and ( w6099 , w6098 , w59 );
and ( w6100 , w6099 , w1244 );
not ( w6101 , w6083 );
and ( w6102 , w6101 , w6100 );
and ( w6103 , w6102 , g11 );
nor ( w6104 , w6072 , w6103 );
and ( w6105 , w6104 , g12 );
and ( w6106 , w6105 , g10 );
and ( w6107 , w6106 , w8765 );
and ( w6108 , w6107 , w8767 );
nor ( w6109 , w6108 , g1 );
and ( w6110 , w6109 , w8845 );
not ( w6111 , w6110 );
and ( w6112 , w6111 , g16 );
not ( w6113 , w6112 );
and ( w6114 , w6113 , w6004 );
and ( w6115 , w4873 , w8767 );
nor ( w6116 , w6115 , g8 );
and ( w6117 , w6116 , w8765 );
not ( w6118 , w6117 );
and ( w6119 , w6118 , w1248 );
not ( w6120 , w6119 );
and ( w6121 , w6120 , g10 );
nor ( w6122 , w6121 , g3 );
and ( w6123 , w6122 , w6062 );
and ( w6124 , w6114 , w6123 );
and ( w6125 , w6124 , w59 );
and ( w6126 , w6125 , w1244 );
not ( w6127 , w6126 );
and ( w6128 , w6127 , g11 );
nor ( w6129 , w5802 , g3 );
and ( w6130 , w6129 , g7 );
and ( w6131 , w3189 , w8767 );
nor ( w6132 , w6131 , g7 );
not ( w6133 , w6132 );
and ( w6134 , w6133 , w17 );
nor ( w6135 , w6134 , g9 );
nor ( w6136 , w6135 , g1 );
nor ( w6137 , w6136 , g8 );
and ( w6138 , w6137 , w8769 );
nor ( w6139 , w6138 , g5 );
and ( w6140 , w6139 , w8742 );
and ( w6141 , w6140 , w408 );
nor ( w6142 , w6141 , g9 );
nor ( w6143 , w6142 , g10 );
and ( w6144 , w6143 , w8767 );
nor ( w6145 , w6144 , g10 );
and ( w6146 , w6145 , w8767 );
nor ( w6147 , w5794 , w6146 );
and ( w6148 , w6085 , w8730 );
and ( w6149 , w6148 , w361 );
nor ( w6150 , w6149 , g8 );
not ( w6151 , w33 );
and ( w6152 , w6150 , w6151 );
and ( w6153 , w6152 , w8765 );
nor ( w6154 , w6153 , g4 );
and ( w6155 , w6154 , w8845 );
and ( w6156 , w6155 , w6030 );
and ( w6157 , w6156 , w8792 );
and ( w6158 , w6147 , w6157 );
and ( w6159 , w6158 , w59 );
not ( w6160 , w5802 );
and ( w6161 , w6159 , w6160 );
not ( w6162 , w6161 );
and ( w6163 , w6162 , g16 );
not ( w6164 , w6163 );
and ( w6165 , w6164 , w6030 );
nor ( w6166 , w6165 , g11 );
nor ( w6167 , w6166 , g3 );
not ( w6168 , w6167 );
and ( w6169 , w6168 , g13 );
nor ( w6170 , w6169 , g1 );
and ( w6171 , w6170 , w8845 );
and ( w6172 , w6171 , w7783 );
nor ( w6173 , w6130 , w6172 );
and ( w6174 , w6173 , g16 );
not ( w6175 , w6174 );
and ( w6176 , w6175 , w6030 );
nor ( w6177 , w6176 , g11 );
nor ( w6178 , w6177 , g3 );
not ( w6179 , w6178 );
and ( w6180 , w6179 , g13 );
nor ( w6181 , w6180 , g1 );
and ( w6182 , w6181 , w8845 );
and ( w6183 , w6182 , w7783 );
and ( w6184 , w6183 , w8735 );
and ( w6185 , w1610 , w8742 );
and ( w6186 , w6184 , w6366 );
not ( w6187 , w6128 );
and ( w6188 , w6187 , w6186 );
not ( w6189 , w6188 );
and ( w6190 , w6189 , g13 );
nor ( w6191 , w6190 , g1 );
and ( w6192 , w6191 , w7783 );
and ( w6193 , w6192 , w8845 );
and ( w6194 , w6193 , w6366 );
nor ( w6195 , w6063 , w6194 );
not ( w6196 , w6195 );
and ( w6197 , w6196 , w6186 );
not ( w6198 , w6060 );
and ( w6199 , w6198 , w6197 );
and ( w6200 , w1429 , w33 );
and ( w6201 , w6200 , w8767 );
nor ( w6202 , w6201 , g9 );
and ( w6203 , w6202 , w8767 );
nor ( w6204 , w6203 , g6 );
and ( w6205 , w6199 , w6204 );
and ( w6206 , w6105 , w8742 );
and ( w6207 , w6206 , w8765 );
and ( w6208 , w6207 , w8767 );
not ( w6209 , w6208 );
and ( w6210 , w6205 , w6209 );
and ( w6211 , w6210 , w1248 );
and ( w6212 , w6197 , w8730 );
not ( w6213 , w6212 );
and ( w6214 , w6213 , g13 );
nor ( w6215 , w6214 , g1 );
and ( w6216 , w6215 , w7783 );
and ( w6217 , w6216 , w8845 );
and ( w6218 , w6217 , w6366 );
nor ( w6219 , w6211 , w6218 );
not ( w6220 , w6219 );
and ( w6221 , w6220 , w27 );
not ( w6222 , w6221 );
and ( w6223 , w6222 , w213 );
nor ( w6224 , w6223 , g1 );
and ( w6225 , w6224 , w7783 );
and ( w6226 , w6225 , w8845 );
not ( w6227 , w6226 );
and ( w6228 , w6227 , g16 );
and ( w6229 , w6197 , w6021 );
not ( w6230 , w6229 );
and ( w6231 , w6230 , g13 );
nor ( w6232 , w6231 , g1 );
and ( w6233 , w6232 , w7783 );
and ( w6234 , w6233 , w8845 );
and ( w6235 , w6234 , w6366 );
not ( w6236 , w6228 );
and ( w6237 , w6236 , w6235 );
and ( w6238 , w6237 , w6021 );
not ( w6239 , w6238 );
and ( w6240 , w6239 , g11 );
not ( w6241 , w6240 );
and ( w6242 , w6241 , w6186 );
not ( w6243 , w6242 );
and ( w6244 , w6243 , g13 );
nor ( w6245 , w6244 , g1 );
and ( w6246 , w6245 , w7783 );
and ( w6247 , w6246 , w8845 );
and ( w6248 , w6247 , w6366 );
and ( w6249 , w8735 , w6248 );
nor ( w6250 , w241 , w6249 );
not ( w6251 , w6250 );
and ( w6252 , w6251 , w17 );
and ( w6253 , w6252 , w8735 );
nor ( w6254 , w6054 , w6253 );
and ( w6255 , w43 , w8742 );
and ( w6256 , w6255 , g3 );
nor ( w6257 , w6256 , w5921 );
nor ( w6258 , w3200 , g6 );
nor ( w6259 , w6258 , g4 );
not ( w6260 , w6259 );
and ( w6261 , w6260 , w471 );
and ( w6262 , w1588 , w1844 );
and ( w6263 , w6262 , w59 );
nor ( w6264 , w6263 , g7 );
and ( w6265 , w6264 , w8860 );
and ( w6266 , w6265 , w8769 );
not ( w6267 , w6266 );
and ( w6268 , w6261 , w6267 );
and ( w6269 , w6268 , g3 );
and ( w6270 , w6269 , w7783 );
not ( w6271 , w6257 );
and ( w6272 , w6271 , w6270 );
and ( w6273 , w7890 , w408 );
and ( w6274 , w6273 , g7 );
and ( w6275 , w240 , w8735 );
and ( w6276 , w6273 , w8767 );
and ( w6277 , w6276 , w8742 );
nor ( w6278 , w6277 , g8 );
not ( w6279 , w6278 );
and ( w6280 , w6279 , g10 );
and ( w6281 , w6280 , w8769 );
and ( w6282 , w6273 , w8735 );
and ( w6283 , w6281 , w6282 );
and ( w6284 , w6275 , w6283 );
and ( w6285 , w6284 , w59 );
nor ( w6286 , w6274 , w6285 );
nor ( w6287 , w6286 , g4 );
and ( w6288 , w6287 , w8845 );
and ( w6289 , w6074 , g12 );
and ( w6290 , w6289 , w8837 );
and ( w6291 , w6290 , w8828 );
not ( w6292 , w6291 );
and ( w6293 , w6292 , w213 );
and ( w6294 , w6293 , g12 );
and ( w6295 , w6294 , w8742 );
and ( w6296 , w6295 , g8 );
and ( w6297 , w6296 , w8819 );
not ( w6298 , w6297 );
and ( w6299 , w6288 , w6298 );
and ( w6300 , w472 , g7 );
and ( w6301 , w6300 , w1260 );
and ( w6302 , w6301 , w8828 );
nor ( w6303 , w6302 , g14 );
and ( w6304 , w6303 , w8765 );
and ( w6305 , w6304 , w8860 );
and ( w6306 , w6305 , w8728 );
and ( w6307 , w6306 , g7 );
nor ( w6308 , w6307 , g6 );
nor ( w6309 , w6308 , g11 );
and ( w6310 , w6309 , w8819 );
nor ( w6311 , w6310 , g1 );
and ( w6312 , w6311 , w8845 );
and ( w6313 , w6299 , w6312 );
and ( w6314 , w6313 , w17 );
and ( w6315 , w6314 , g10 );
nor ( w6316 , w6315 , g11 );
and ( w6317 , w6316 , w8828 );
nor ( w6318 , w6317 , g1 );
and ( w6319 , w6318 , w8845 );
nor ( w6320 , w6272 , w6319 );
not ( w6321 , w6320 );
and ( w6322 , w6321 , g10 );
and ( w6323 , w3559 , w8767 );
not ( w6324 , w6323 );
and ( w6325 , w6324 , g9 );
and ( w6326 , w6325 , w8767 );
and ( w6327 , w6335 , g9 );
and ( w6328 , w40 , g3 );
and ( w6329 , w6328 , w8765 );
nor ( w6330 , w6327 , w6329 );
nor ( w6331 , w6330 , g4 );
and ( w6332 , w6331 , w2687 );
and ( w6333 , w6332 , w8742 );
and ( w6334 , w6333 , w8845 );
not ( w6335 , w6326 );
and ( w6336 , w6335 , g3 );
and ( w6337 , w6334 , w6336 );
and ( w6338 , w6336 , g7 );
nor ( w6339 , w6337 , w6338 );
and ( w6340 , w3559 , g9 );
nor ( w6341 , w6340 , w6270 );
nor ( w6342 , w6341 , g10 );
and ( w6343 , w6342 , w8845 );
and ( w6344 , w6343 , w7783 );
not ( w6345 , w6339 );
and ( w6346 , w6345 , w6344 );
and ( w6347 , w1575 , w1579 );
not ( w6348 , w6347 );
and ( w6349 , w6348 , g18 );
and ( w6350 , w6349 , g9 );
and ( w6351 , w6350 , w8767 );
nor ( w6352 , w6351 , g10 );
and ( w6353 , w6352 , w3200 );
and ( w6354 , w6353 , w7783 );
and ( w6355 , w8792 , w6354 );
nor ( w6356 , w6346 , w6355 );
and ( w6357 , w6630 , g11 );
not ( w6358 , w6357 );
and ( w6359 , w6358 , w5803 );
and ( w6360 , w6359 , g3 );
nor ( w6361 , w6360 , w6248 );
and ( w6362 , w6361 , g13 );
nor ( w6363 , w6362 , g1 );
and ( w6364 , w6363 , w7783 );
and ( w6365 , w6364 , w8845 );
not ( w6366 , w6185 );
and ( w6367 , w6365 , w6366 );
not ( w6368 , w6356 );
and ( w6369 , w6368 , w6367 );
nor ( w6370 , w6322 , w6369 );
nor ( w6371 , w6370 , g2 );
nor ( w6372 , w6371 , g16 );
not ( w6373 , w6372 );
and ( w6374 , w6373 , w6367 );
nor ( w6375 , g9 , w6374 );
not ( w6376 , w6375 );
and ( w6377 , w6376 , g10 );
nor ( w6378 , w6377 , w6369 );
not ( w6379 , w6378 );
and ( w6380 , w6379 , w6367 );
nor ( w6381 , w1786 , w6380 );
and ( w6382 , w6381 , w7783 );
nor ( w6383 , w6382 , g6 );
and ( w6384 , w6383 , w8735 );
and ( w6385 , w6384 , w8792 );
not ( w6386 , w6254 );
and ( w6387 , w6386 , w6385 );
and ( w6388 , w6387 , w27 );
and ( w6389 , w471 , w8742 );
and ( w6390 , w6389 , g8 );
and ( w6391 , w6390 , g2 );
and ( w6392 , w6391 , w8769 );
and ( w6393 , w6392 , g10 );
and ( w6394 , w6393 , w8860 );
nor ( w6395 , w6394 , g5 );
and ( w6396 , w6395 , w8860 );
and ( w6397 , w6396 , w8742 );
and ( w6398 , w6397 , g8 );
and ( w6399 , w1982 , w8735 );
and ( w6400 , w6399 , w8765 );
not ( w6401 , w6398 );
and ( w6402 , w6401 , w6400 );
and ( w6403 , w6402 , g2 );
and ( w6404 , w7783 , g7 );
and ( w6405 , w6404 , w8735 );
not ( w6406 , w6303 );
and ( w6407 , w6406 , w6405 );
not ( w6408 , w6407 );
and ( w6409 , w6408 , g7 );
nor ( w6410 , w6409 , g9 );
and ( w6411 , w6410 , w8860 );
nor ( w6412 , w6411 , g12 );
and ( w6413 , w6412 , w8837 );
and ( w6414 , w6413 , w8819 );
nor ( w6415 , w6414 , g1 );
and ( w6416 , w6415 , w8845 );
and ( w6417 , w6416 , w8735 );
nor ( w6418 , g3 , w6417 );
and ( w6419 , w6418 , w8765 );
and ( w6420 , w6419 , w8728 );
not ( w6421 , w6420 );
and ( w6422 , w6421 , w6380 );
nor ( w6423 , w6422 , g16 );
not ( w6424 , w6423 );
and ( w6425 , w6424 , w6367 );
and ( w6426 , w6425 , w8769 );
and ( w6427 , w6426 , w8860 );
nor ( w6428 , w6427 , g5 );
and ( w6429 , w6428 , w8860 );
nor ( w6430 , w6429 , g7 );
nor ( w6431 , w6430 , g7 );
not ( w6432 , w6431 );
and ( w6433 , w6432 , g8 );
not ( w6434 , w6433 );
and ( w6435 , w6434 , g8 );
not ( w6436 , w5098 );
and ( w6437 , w6436 , w27 );
nor ( w6438 , w6437 , g4 );
not ( w6439 , w6438 );
and ( w6440 , w6439 , w5819 );
and ( w6441 , w6440 , w8735 );
not ( w6442 , w6435 );
and ( w6443 , w6442 , w6441 );
and ( w6444 , w6443 , w8845 );
and ( w6445 , w6444 , w8792 );
nor ( w6446 , w6403 , w6445 );
not ( w6447 , w6446 );
and ( w6448 , w6447 , g10 );
and ( w6449 , w6448 , w33 );
and ( w6450 , w6449 , w8845 );
nor ( w6451 , w1347 , w5891 );
nor ( w6452 , w6451 , g3 );
nor ( w6453 , w6452 , g16 );
not ( w6454 , w6453 );
and ( w6455 , w6454 , w33 );
nor ( w6456 , g4 , w6367 );
and ( w6457 , w6456 , w7783 );
and ( w6458 , w6457 , w8769 );
and ( w6459 , w6455 , w6519 );
not ( w6460 , w6459 );
and ( w6461 , w6460 , g11 );
and ( w6462 , w6461 , g13 );
nor ( w6463 , w6462 , g6 );
and ( w6464 , w6463 , w8735 );
and ( w6465 , w6464 , w8792 );
nor ( w6466 , w6465 , w1408 );
and ( w6467 , w27 , g10 );
and ( w6468 , w6467 , w59 );
nor ( w6469 , w6468 , g7 );
and ( w6470 , w6469 , w8860 );
not ( w6471 , w6470 );
and ( w6472 , w6471 , g10 );
and ( w6473 , w3408 , w8860 );
not ( w6474 , w6473 );
and ( w6475 , w6472 , w6474 );
not ( w6476 , w6475 );
and ( w6477 , w6476 , g11 );
and ( w6478 , w6477 , g13 );
and ( w6479 , w6478 , g12 );
nor ( w6480 , w6479 , g3 );
nor ( w6481 , w2075 , w6480 );
nor ( w6482 , w6481 , g1 );
and ( w6483 , w6482 , w400 );
nor ( w6484 , w1248 , g5 );
nor ( w6485 , w1609 , w6484 );
not ( w6486 , w1235 );
and ( w6487 , w6485 , w6486 );
and ( w6488 , w6487 , w7783 );
and ( w6489 , w6488 , w8792 );
and ( w6490 , w6489 , w6021 );
nor ( w6491 , w6490 , w6367 );
not ( w6492 , w6491 );
and ( w6493 , w6492 , w1260 );
and ( w6494 , w6493 , g10 );
nor ( w6495 , w6483 , w6494 );
not ( w6496 , w6495 );
and ( w6497 , w6496 , g10 );
not ( w6498 , w6497 );
and ( w6499 , w6498 , g10 );
and ( w6500 , w6499 , g16 );
not ( w6501 , w6500 );
and ( w6502 , w6501 , w5902 );
not ( w6503 , w6502 );
and ( w6504 , w6503 , w213 );
nor ( w6505 , w6504 , w6458 );
not ( w6506 , w6505 );
and ( w6507 , w6506 , g11 );
and ( w6508 , w6507 , g13 );
and ( w6509 , w6508 , g12 );
nor ( w6510 , w6509 , g6 );
and ( w6511 , w6510 , w8735 );
and ( w6512 , w6511 , w8792 );
not ( w6513 , w6466 );
and ( w6514 , w6513 , w6512 );
not ( w6515 , w6514 );
and ( w6516 , w6515 , w213 );
not ( w6517 , w6516 );
and ( w6518 , w6517 , w6275 );
not ( w6519 , w6458 );
and ( w6520 , w6518 , w6519 );
not ( w6521 , w6520 );
and ( w6522 , w6521 , g11 );
nor ( w6523 , w33 , w1408 );
not ( w6524 , w6523 );
and ( w6525 , w6524 , g2 );
nor ( w6526 , w6525 , w5819 );
nor ( w6527 , w6526 , g9 );
not ( w6528 , w5803 );
and ( w6529 , g10 , w6528 );
and ( w6530 , w6529 , w7783 );
nor ( w6531 , w6530 , g3 );
and ( w6532 , w6531 , g7 );
nor ( w6533 , g10 , g6 );
and ( w6534 , w7890 , w6533 );
and ( w6535 , w6534 , w8767 );
nor ( w6536 , w6535 , g10 );
nor ( w6537 , w6536 , g8 );
nor ( w6538 , w6537 , g8 );
nor ( w6539 , w6538 , g1 );
and ( w6540 , w1367 , w8860 );
and ( w6541 , w6540 , w8769 );
not ( w6542 , w6541 );
and ( w6543 , w6539 , w6542 );
not ( w6544 , w6543 );
and ( w6545 , w6544 , w213 );
not ( w6546 , w5876 );
and ( w6547 , w6545 , w6546 );
not ( w6548 , w6547 );
and ( w6549 , w6548 , g2 );
and ( w6550 , w6549 , w400 );
nor ( w6551 , w6159 , g5 );
and ( w6552 , w6551 , w8860 );
nor ( w6553 , w6552 , w5802 );
and ( w6554 , w6553 , w7783 );
nor ( w6555 , w6554 , g11 );
and ( w6556 , w6555 , g13 );
nor ( w6557 , w6556 , g6 );
and ( w6558 , w6557 , w8735 );
and ( w6559 , w6558 , w8792 );
nor ( w6560 , w6550 , w6559 );
nor ( w6561 , w6560 , g7 );
not ( w6562 , w6561 );
and ( w6563 , w6562 , g16 );
and ( w6564 , w6563 , w8837 );
and ( w6565 , w6564 , g13 );
and ( w6566 , w6565 , g12 );
nor ( w6567 , w6566 , g6 );
and ( w6568 , w6567 , w8735 );
and ( w6569 , w6568 , w8792 );
nor ( w6570 , w6532 , w6569 );
and ( w6571 , w6570 , w8837 );
and ( w6572 , w6571 , g13 );
and ( w6573 , w6572 , g12 );
nor ( w6574 , w6573 , g6 );
and ( w6575 , w6574 , w8735 );
and ( w6576 , w6575 , w8792 );
and ( w6577 , w6527 , w6576 );
not ( w6578 , w6522 );
and ( w6579 , w6578 , w6577 );
not ( w6580 , w6579 );
and ( w6581 , w6580 , g13 );
and ( w6582 , w6581 , g12 );
nor ( w6583 , w6582 , g6 );
and ( w6584 , w6583 , w361 );
and ( w6585 , w6584 , w408 );
and ( w6586 , w6450 , w6585 );
not ( w6587 , w4418 );
and ( w6588 , w6587 , g4 );
nor ( w6589 , w6588 , g9 );
and ( w6590 , w6589 , w8845 );
and ( w6591 , w6590 , w8792 );
and ( w6592 , w6591 , w5800 );
not ( w6593 , w6592 );
and ( w6594 , w6593 , g2 );
nor ( w6595 , w6594 , g10 );
and ( w6596 , w6595 , w6585 );
nor ( w6597 , w6586 , w6596 );
not ( w6598 , w6597 );
and ( w6599 , w6388 , w6598 );
not ( w6600 , w6599 );
and ( w6601 , w6046 , w6600 );
nor ( w6602 , w6601 , w6597 );
not ( w6603 , w6041 );
and ( w6604 , w6603 , w6602 );
not ( w6605 , w5905 );
and ( w6606 , w6605 , w6604 );
not ( w6607 , w5838 );
and ( w6608 , w6607 , w6606 );
nor ( w6609 , w6608 , g13 );
not ( w6610 , w6609 );
and ( w6611 , w6610 , w6606 );
nor ( w6612 , w6611 , g16 );
nor ( w6613 , w6612 , g3 );
nor ( w6614 , w6613 , g12 );
not ( w6615 , w6614 );
and ( w6616 , w6615 , w6602 );
not ( w6617 , w5828 );
and ( w6618 , w6617 , w6616 );
nor ( w6619 , w5738 , w6618 );
nor ( w6620 , w6619 , g6 );
and ( w6621 , w6620 , g2 );
and ( w6622 , w6621 , w8792 );
nor ( w6623 , w5746 , w6622 );
and ( w6624 , w2585 , w8767 );
not ( w6625 , w6624 );
and ( w6626 , w6625 , w1366 );
not ( w6627 , w6626 );
and ( w6628 , w6627 , w4793 );
and ( w6629 , w1353 , w8845 );
not ( w6630 , w5891 );
and ( w6631 , w6630 , g13 );
nor ( w6632 , w6631 , g1 );
nor ( w6633 , w4357 , w6632 );
and ( w6634 , w1516 , g10 );
and ( w6635 , w8765 , w2585 );
and ( w6636 , w6635 , w8730 );
nor ( w6637 , w1408 , g10 );
nor ( w6638 , g2 , w6637 );
and ( w6639 , w6638 , g6 );
and ( w6640 , w6639 , w8792 );
not ( w6641 , w1366 );
and ( w6642 , g2 , w6641 );
not ( w6643 , w6642 );
and ( w6644 , w6643 , w2669 );
and ( w6645 , w4359 , w8730 );
not ( w6646 , w6644 );
and ( w6647 , w6646 , w6645 );
and ( w6648 , w6647 , w1408 );
not ( w6649 , w6648 );
and ( w6650 , w6649 , g11 );
nor ( w6651 , w6650 , g9 );
nor ( w6652 , w1347 , w6651 );
and ( w6653 , w243 , g3 );
and ( w6654 , w6653 , w8742 );
and ( w6655 , w6654 , w59 );
nor ( w6656 , w6655 , g7 );
not ( w6657 , w6656 );
and ( w6658 , w6657 , g10 );
and ( w6659 , w6658 , w33 );
nor ( w6660 , w6659 , g4 );
and ( w6661 , w6660 , w8769 );
and ( w6662 , w6661 , g10 );
nor ( w6663 , w6662 , g6 );
and ( w6664 , w6663 , g2 );
and ( w6665 , w6631 , w8828 );
nor ( w6666 , w6665 , g1 );
nor ( w6667 , w6664 , w6666 );
not ( w6668 , w6618 );
and ( w6669 , w6667 , w6668 );
nor ( w6670 , w6669 , g6 );
not ( w6671 , w6670 );
and ( w6672 , w6671 , g11 );
nor ( w6673 , w5149 , w2224 );
not ( w6674 , w6673 );
and ( w6675 , w6674 , g2 );
nor ( w6676 , w4416 , w104 );
nor ( w6677 , w6676 , g2 );
and ( w6678 , w6677 , w8765 );
not ( w6679 , w6588 );
and ( w6680 , w6679 , g6 );
nor ( w6681 , w2844 , w6618 );
nor ( w6682 , w6681 , g3 );
and ( w6683 , w6682 , w8730 );
and ( w6684 , w6683 , w8765 );
and ( w6685 , w6684 , w8792 );
and ( w6686 , w6680 , w6685 );
nor ( w6687 , w6686 , w6618 );
not ( w6688 , w5767 );
and ( w6689 , w6687 , w6688 );
nor ( w6690 , w6689 , g10 );
and ( w6691 , w6690 , w8765 );
nor ( w6692 , w6691 , g9 );
not ( w6693 , w6692 );
and ( w6694 , w6693 , w1588 );
and ( w6695 , w6694 , w8730 );
nor ( w6696 , w6695 , g10 );
nor ( w6697 , g3 , w291 );
nor ( w6698 , w6697 , g9 );
nor ( w6699 , w6698 , g4 );
not ( w6700 , w6699 );
and ( w6701 , w6700 , g2 );
and ( w6702 , w6701 , g7 );
not ( w6703 , w6702 );
and ( w6704 , w6703 , g2 );
and ( w6705 , w6704 , g7 );
not ( w6706 , w6705 );
and ( w6707 , w6706 , g6 );
nor ( w6708 , w4900 , g6 );
and ( w6709 , w6708 , g3 );
nor ( w6710 , w6709 , w6618 );
nor ( w6711 , w6710 , g9 );
and ( w6712 , w6711 , w8792 );
nor ( w6713 , w6707 , w6712 );
nor ( w6714 , w6713 , g1 );
and ( w6715 , w6714 , g10 );
nor ( w6716 , g4 , w291 );
not ( w6717 , w6716 );
and ( w6718 , w6717 , g2 );
and ( w6719 , w6718 , w8792 );
and ( w6720 , w6719 , g10 );
nor ( w6721 , w1898 , w291 );
nor ( w6722 , w6721 , g10 );
and ( w6723 , w6722 , g2 );
and ( w6724 , w6723 , w8792 );
and ( w6725 , w6724 , w408 );
nor ( w6726 , w6720 , w6725 );
nor ( w6727 , w6726 , g3 );
and ( w6728 , w6727 , w408 );
and ( w6729 , w6728 , w8742 );
and ( w6730 , w6729 , w8730 );
and ( w6731 , w6730 , g4 );
nor ( w6732 , w6731 , g3 );
and ( w6733 , w6732 , g4 );
and ( w6734 , w6733 , g2 );
not ( w6735 , w6734 );
and ( w6736 , w6735 , g5 );
and ( w6737 , w6736 , g6 );
and ( w6738 , w6737 , w8742 );
and ( w6739 , w6738 , w8765 );
nor ( w6740 , w6739 , g7 );
and ( w6741 , w6740 , g5 );
not ( w6742 , w6741 );
and ( w6743 , w6742 , w6714 );
and ( w6744 , w6743 , g6 );
nor ( w6745 , w6744 , w6712 );
not ( w6746 , w6715 );
and ( w6747 , w6746 , w6745 );
and ( w6748 , w3024 , w408 );
and ( w6749 , w6748 , w8792 );
not ( w6750 , w6747 );
and ( w6751 , w6750 , w6749 );
nor ( w6752 , w6751 , g9 );
nor ( w6753 , w6752 , g1 );
and ( w6754 , w6753 , g10 );
not ( w6755 , w4793 );
and ( w6756 , w6755 , g13 );
and ( w6757 , w6756 , w8828 );
nor ( w6758 , w6757 , g1 );
nor ( w6759 , w6754 , w6758 );
nor ( w6760 , w6696 , w6759 );
and ( w6761 , w6678 , w6760 );
nor ( w6762 , w6675 , w6761 );
and ( w6763 , w6762 , w8837 );
nor ( w6764 , w6763 , g9 );
not ( w6765 , w6764 );
and ( w6766 , w6765 , w213 );
not ( w6767 , w6766 );
and ( w6768 , w6767 , w6760 );
not ( w6769 , w6768 );
and ( w6770 , w6769 , g13 );
and ( w6771 , w6770 , w8828 );
nor ( w6772 , w6771 , g1 );
not ( w6773 , w6672 );
and ( w6774 , w6773 , w6772 );
and ( w6775 , w6774 , w8765 );
not ( w6776 , w6775 );
and ( w6777 , w6776 , w213 );
not ( w6778 , w6777 );
and ( w6779 , w6778 , w6760 );
not ( w6780 , w6779 );
and ( w6781 , w6780 , g13 );
and ( w6782 , w6781 , w8828 );
nor ( w6783 , w6782 , g1 );
not ( w6784 , w6652 );
and ( w6785 , w6784 , w6783 );
and ( w6786 , w6533 , w8767 );
and ( w6787 , w6786 , w8735 );
nor ( w6788 , w6787 , g8 );
and ( w6789 , w6788 , w8735 );
nor ( w6790 , g10 , w6789 );
and ( w6791 , w6790 , w8845 );
and ( w6792 , w6791 , w8730 );
and ( w6793 , w6792 , w8845 );
and ( w6794 , w3470 , w6793 );
and ( w6795 , w6794 , g11 );
and ( w6796 , w6795 , g9 );
and ( w6797 , w6796 , g2 );
and ( w6798 , w6797 , g17 );
and ( w6799 , w6798 , g15 );
and ( w6800 , w6799 , g16 );
and ( w6801 , w6800 , g14 );
not ( w6802 , w6801 );
and ( w6803 , w6802 , g13 );
not ( w6804 , w6803 );
and ( w6805 , w6804 , w400 );
and ( w6806 , w6805 , w8792 );
nor ( w6807 , w6785 , w6806 );
not ( w6808 , w6807 );
and ( w6809 , w6808 , g2 );
nor ( w6810 , w6809 , w6666 );
not ( w6811 , w6810 );
and ( w6812 , w6811 , g3 );
nor ( w6813 , w6812 , w6618 );
nor ( w6814 , w6813 , g6 );
not ( w6815 , w6814 );
and ( w6816 , w6815 , g11 );
not ( w6817 , w6816 );
and ( w6818 , w6817 , w6772 );
and ( w6819 , w6818 , w8765 );
not ( w6820 , w6819 );
and ( w6821 , w6820 , w213 );
not ( w6822 , w6821 );
and ( w6823 , w6822 , w6760 );
not ( w6824 , w6823 );
and ( w6825 , w6824 , g13 );
and ( w6826 , w6825 , w8828 );
nor ( w6827 , w6826 , g1 );
nor ( w6828 , w6640 , w6827 );
not ( w6829 , w6828 );
and ( w6830 , w6829 , w6772 );
and ( w6831 , w6830 , w8765 );
and ( w6832 , w6831 , w6760 );
nor ( w6833 , w6636 , w6832 );
not ( w6834 , w6833 );
and ( w6835 , w6834 , g6 );
nor ( w6836 , w6835 , w6827 );
and ( w6837 , w6836 , g11 );
not ( w6838 , w6837 );
and ( w6839 , w6838 , w6772 );
nor ( w6840 , w3337 , w6839 );
not ( w6841 , w6840 );
and ( w6842 , w6841 , w6760 );
nor ( w6843 , w6634 , w6842 );
not ( w6844 , w6843 );
and ( w6845 , w6844 , g10 );
nor ( w6846 , w6328 , w1552 );
nor ( w6847 , w6846 , g10 );
and ( w6848 , w6847 , w7783 );
not ( w6849 , w6848 );
and ( w6850 , w6849 , g11 );
not ( w6851 , w1589 );
and ( w6852 , w6851 , g3 );
not ( w6853 , w6852 );
and ( w6854 , w6853 , g9 );
nor ( w6855 , w6854 , w6839 );
not ( w6856 , w6855 );
and ( w6857 , w6856 , w6760 );
not ( w6858 , w6850 );
and ( w6859 , w6858 , w6857 );
and ( w6860 , w6859 , g9 );
nor ( w6861 , w6860 , w6839 );
not ( w6862 , w6845 );
and ( w6863 , w6862 , w6861 );
nor ( w6864 , w6863 , g2 );
not ( w6865 , w6633 );
and ( w6866 , w6865 , w6864 );
and ( w6867 , w6866 , g10 );
not ( w6868 , w6867 );
and ( w6869 , w6868 , w6861 );
not ( w6870 , w6629 );
and ( w6871 , w6870 , w6869 );
not ( w6872 , w6871 );
and ( w6873 , w6872 , w6857 );
nor ( w6874 , w1517 , w6873 );
nor ( w6875 , w6874 , g10 );
and ( w6876 , w6875 , g2 );
not ( w6877 , w6876 );
and ( w6878 , w6877 , w6869 );
not ( w6879 , w6878 );
and ( w6880 , w6879 , w6857 );
and ( w6881 , w6628 , w6880 );
and ( w6882 , w6881 , g2 );
not ( w6883 , w6882 );
and ( w6884 , w6883 , w6869 );
and ( w6885 , w8374 , w6884 );
nor ( w6886 , w6623 , w6885 );
and ( w6887 , w6886 , w8765 );
and ( w6888 , w6887 , w8860 );
nor ( w6889 , w5737 , w6888 );
and ( w6890 , g4 , w8765 );
and ( w6891 , w6890 , g3 );
nor ( w6892 , w6891 , w6618 );
nor ( w6893 , w6892 , g6 );
nor ( w6894 , w6893 , g6 );
not ( w6895 , w1845 );
and ( w6896 , w6894 , w6895 );
not ( w6897 , w6896 );
and ( w6898 , w6897 , g2 );
and ( w6899 , w6898 , w6972 );
not ( w6900 , w6889 );
and ( w6901 , w6900 , w6899 );
nor ( w6902 , w6901 , g9 );
not ( w6903 , w6902 );
and ( w6904 , w6903 , g2 );
and ( w6905 , w6904 , w6972 );
nor ( w6906 , w5375 , g3 );
not ( w6907 , w6906 );
and ( w6908 , w6907 , w17 );
nor ( w6909 , w6908 , g5 );
and ( w6910 , w6909 , w8742 );
and ( w6911 , w6910 , w8860 );
nor ( w6912 , w6911 , g1 );
and ( w6913 , w6912 , w8765 );
and ( w6914 , w6913 , g3 );
not ( w6915 , w6914 );
and ( w6916 , w6915 , g3 );
not ( w6917 , w6916 );
and ( w6918 , w6917 , g6 );
and ( w6919 , w6711 , w6972 );
nor ( w6920 , w6918 , w6919 );
nor ( w6921 , g6 , w6919 );
nor ( w6922 , w6921 , w6885 );
not ( w6923 , w6920 );
and ( w6924 , w6923 , w6922 );
and ( w6925 , w6924 , w8765 );
and ( w6926 , w6925 , g2 );
nor ( w6927 , g6 , w6711 );
nor ( w6928 , w6927 , g9 );
and ( w6929 , w6928 , w4833 );
and ( w6930 , w6632 , g3 );
nor ( w6931 , w6930 , w6618 );
nor ( w6932 , w6931 , w6458 );
and ( w6933 , w6932 , w8845 );
not ( w6934 , w6933 );
and ( w6935 , w6934 , g11 );
nor ( w6936 , w6935 , g2 );
and ( w6937 , w6936 , w8765 );
and ( w6938 , w6929 , w6937 );
and ( w6939 , w5803 , w6938 );
nor ( w6940 , g6 , w6939 );
and ( w6941 , w6940 , g16 );
nor ( w6942 , w6941 , w6885 );
and ( w6943 , w6942 , w7783 );
and ( w6944 , w6943 , w8765 );
nor ( w6945 , g1 , w6944 );
nor ( w6946 , w6945 , g2 );
not ( w6947 , w3683 );
and ( w6948 , w6947 , g13 );
and ( w6949 , w6948 , w8845 );
and ( w6950 , w6949 , w8828 );
nor ( w6951 , w6950 , g15 );
and ( w6952 , w6951 , g1 );
and ( w6953 , w41 , w6972 );
and ( w6954 , w4570 , w7783 );
and ( w6955 , w6954 , w59 );
nor ( w6956 , w6955 , g7 );
and ( w6957 , w6956 , w8860 );
and ( w6958 , w6957 , w8769 );
not ( w6959 , w6958 );
and ( w6960 , w6959 , g6 );
and ( w6961 , w6960 , w526 );
and ( w6962 , w6961 , w1489 );
and ( w6963 , w6944 , g3 );
not ( w6964 , w6963 );
and ( w6965 , w6964 , g13 );
not ( w6966 , w6965 );
and ( w6967 , w6966 , g3 );
and ( w6968 , w6967 , w7783 );
nor ( w6969 , w6968 , g12 );
and ( w6970 , w3736 , w6944 );
and ( w6971 , w7783 , g3 );
not ( w6972 , w6885 );
and ( w6973 , w6971 , w6972 );
and ( w6974 , w520 , w6973 );
nor ( w6975 , w516 , w6618 );
not ( w6976 , w6975 );
and ( w6977 , w6976 , w2190 );
and ( w6978 , w6977 , w1844 );
nor ( w6979 , w6974 , w6978 );
and ( w6980 , w6979 , g12 );
nor ( w6981 , w6980 , g9 );
nor ( w6982 , w6970 , w6981 );
not ( w6983 , w6926 );
and ( w6984 , w6983 , w6982 );
nor ( w6985 , w6969 , w6984 );
and ( w6986 , w6270 , w6985 );
and ( w6987 , g4 , w41 );
nor ( w6988 , w6987 , w27 );
nor ( w6989 , w6988 , g3 );
nor ( w6990 , g3 , w6618 );
and ( w6991 , w6990 , w8845 );
not ( w6992 , w6991 );
and ( w6993 , w41 , w6992 );
and ( w6994 , w6989 , w6993 );
nor ( w6995 , w6986 , w6994 );
and ( w6996 , w6995 , w8837 );
nor ( w6997 , w6996 , g2 );
and ( w6998 , w6997 , w7006 );
nor ( w6999 , w6962 , w6998 );
not ( w7000 , w6999 );
and ( w7001 , w7000 , w6985 );
and ( w7002 , w7001 , w6971 );
nor ( w7003 , w7002 , w6994 );
and ( w7004 , w7003 , w8837 );
nor ( w7005 , w7004 , g2 );
not ( w7006 , w6984 );
and ( w7007 , w7005 , w7006 );
and ( w7008 , w6953 , w7007 );
nor ( w7009 , w6926 , w7008 );
not ( w7010 , w6952 );
and ( w7011 , w7010 , w7009 );
nor ( w7012 , w7011 , g9 );
and ( w7013 , w6946 , w7012 );
nor ( w7014 , w6926 , w7013 );
and ( w7015 , w1588 , w7014 );
not ( w7016 , w7015 );
and ( w7017 , w7016 , g2 );
nor ( w7018 , w7017 , w7013 );
not ( w7019 , w7018 );
and ( w7020 , w7019 , w7012 );
nor ( w7021 , g9 , w7020 );
nor ( w7022 , w6885 , w7021 );
and ( w7023 , w7022 , w7783 );
and ( w7024 , w7023 , g9 );
nor ( w7025 , w7024 , w7020 );
not ( w7026 , w7025 );
and ( w7027 , w7026 , w1489 );
nor ( w7028 , w6359 , w7020 );
and ( w7029 , w7028 , g13 );
nor ( w7030 , w7029 , w7021 );
not ( w7031 , w7030 );
and ( w7032 , w7031 , g16 );
nor ( w7033 , w7032 , w7021 );
and ( w7034 , w7033 , w8792 );
nor ( w7035 , w7027 , w7034 );
nor ( w7036 , w7035 , g2 );
and ( w7037 , w7036 , w7022 );
nor ( w7038 , w6905 , w7037 );
and ( w7039 , w7038 , w7345 );
and ( w7040 , w7973 , g8 );
not ( w7041 , w7040 );
and ( w7042 , w7039 , w7041 );
and ( w7043 , w8792 , w7038 );
nor ( w7044 , w7043 , w7021 );
and ( w7045 , w7044 , g2 );
and ( w7046 , w7045 , g1 );
not ( w7047 , w7046 );
and ( w7048 , w7047 , w7038 );
not ( w7049 , w7048 );
and ( w7050 , w7049 , g6 );
and ( w7051 , w7050 , g2 );
and ( w7052 , w7051 , g9 );
nor ( w7053 , w7052 , w7020 );
not ( w7054 , w7053 );
and ( w7055 , w7054 , g6 );
and ( w7056 , w7364 , w7055 );
nor ( w7057 , w7056 , g13 );
and ( w7058 , w7044 , w7783 );
and ( w7059 , w7058 , w8730 );
and ( w7060 , w7059 , g3 );
and ( w7061 , w7060 , g9 );
nor ( w7062 , w7061 , w7020 );
not ( w7063 , w7062 );
and ( w7064 , w7063 , g17 );
and ( w7065 , w7064 , w4849 );
not ( w7066 , w7065 );
and ( w7067 , w7066 , w7038 );
and ( w7068 , w7067 , w7039 );
and ( w7069 , w7068 , g16 );
not ( w7070 , w59 );
and ( w7071 , w7039 , w7070 );
nor ( w7072 , w299 , w59 );
and ( w7073 , w7071 , w7072 );
nor ( w7074 , w7043 , g4 );
and ( w7075 , w7074 , g12 );
and ( w7076 , w7075 , w8382 );
and ( w7077 , w7076 , g14 );
and ( w7078 , w7077 , w7044 );
and ( w7079 , w7078 , g3 );
and ( w7080 , w7079 , g9 );
nor ( w7081 , w7080 , w7020 );
not ( w7082 , w7081 );
and ( w7083 , w7082 , g17 );
and ( w7084 , w7083 , w4849 );
not ( w7085 , w7084 );
and ( w7086 , w7085 , w7038 );
and ( w7087 , w7086 , w7039 );
and ( w7088 , w7087 , w8837 );
not ( w7089 , w7088 );
and ( w7090 , w7089 , w2585 );
not ( w7091 , w7090 );
and ( w7092 , w7091 , g6 );
nor ( w7093 , w7092 , w2669 );
not ( w7094 , w7093 );
and ( w7095 , w7094 , w7038 );
and ( w7096 , w7095 , w7345 );
not ( w7097 , w7096 );
and ( w7098 , w7097 , g2 );
and ( w7099 , w2669 , w7038 );
and ( w7100 , w7099 , w7345 );
not ( w7101 , w7100 );
and ( w7102 , w7101 , w104 );
not ( w7103 , w7102 );
and ( w7104 , w7103 , w7039 );
nor ( w7105 , w7104 , g2 );
and ( w7106 , w7105 , w7216 );
nor ( w7107 , w7106 , w7020 );
and ( w7108 , w7107 , w7038 );
and ( w7109 , w7108 , w8828 );
nor ( w7110 , w7109 , w7021 );
and ( w7111 , w7110 , w7044 );
not ( w7112 , w7111 );
and ( w7113 , w7112 , g13 );
not ( w7114 , w7098 );
and ( w7115 , w7114 , w7113 );
and ( w7116 , w7115 , w8828 );
and ( w7117 , w7073 , w7116 );
not ( w7118 , w7117 );
and ( w7119 , w7118 , w7044 );
and ( w7120 , w7044 , w8742 );
and ( w7121 , w7120 , g5 );
and ( w7122 , w7044 , w8769 );
and ( w7123 , w7122 , w1609 );
nor ( w7124 , w7121 , w7123 );
nor ( w7125 , w7124 , g4 );
and ( w7126 , w7125 , g10 );
and ( w7127 , w7126 , g18 );
and ( w7128 , w7127 , g12 );
not ( w7129 , w7128 );
and ( w7130 , w7039 , w7129 );
not ( w7131 , w7130 );
and ( w7132 , w7131 , g3 );
and ( w7133 , w7132 , g9 );
nor ( w7134 , w7133 , w7020 );
not ( w7135 , w7134 );
and ( w7136 , w7135 , g17 );
and ( w7137 , w7136 , w4849 );
not ( w7138 , w7137 );
and ( w7139 , w7138 , w7038 );
and ( w7140 , w7139 , w7039 );
not ( w7141 , g14 );
and ( w7142 , w7140 , w7141 );
and ( w7143 , w8223 , w7044 );
and ( w7144 , w7143 , g17 );
and ( w7145 , w7144 , g12 );
and ( w7146 , w7145 , g3 );
and ( w7147 , w7146 , w8860 );
not ( w7148 , w7147 );
and ( w7149 , w7039 , w7148 );
not ( w7150 , w7149 );
and ( w7151 , w7150 , g10 );
not ( w7152 , w1613 );
and ( w7153 , w7152 , w7038 );
and ( w7154 , w7153 , w7039 );
nor ( w7155 , w7154 , g4 );
and ( w7156 , w7155 , g12 );
nor ( w7157 , w7156 , w7020 );
and ( w7158 , w7157 , w7038 );
not ( w7159 , w7158 );
and ( w7160 , w7159 , w7044 );
and ( w7161 , w7160 , g17 );
nor ( w7162 , w7161 , w7020 );
and ( w7163 , w7162 , w7039 );
not ( w7164 , w7163 );
and ( w7165 , w7164 , w4849 );
not ( w7166 , w7165 );
and ( w7167 , w7166 , w7038 );
and ( w7168 , w7167 , w7039 );
nor ( w7169 , w7168 , g10 );
not ( w7170 , w7169 );
and ( w7171 , w7170 , w7039 );
and ( w7172 , w7171 , g13 );
not ( w7173 , w7151 );
and ( w7174 , w7173 , w7172 );
not ( w7175 , w7174 );
and ( w7176 , w7175 , w7044 );
nor ( w7177 , w7176 , g18 );
and ( w7178 , w7177 , g14 );
nor ( w7179 , w7178 , w7021 );
and ( w7180 , w7179 , w7216 );
and ( w7181 , w7180 , g6 );
not ( w7182 , w7181 );
and ( w7183 , w7182 , g6 );
nor ( w7184 , w7183 , w7021 );
and ( w7185 , w7184 , w7216 );
not ( w7186 , w2669 );
and ( w7187 , w7185 , w7186 );
not ( w7188 , w7187 );
and ( w7189 , w7188 , w7038 );
and ( w7190 , w7189 , w7345 );
and ( w7191 , w7190 , g13 );
nor ( w7192 , w7142 , w7191 );
and ( w7193 , w7192 , g6 );
not ( w7194 , w7193 );
and ( w7195 , w7194 , g6 );
nor ( w7196 , w7195 , w2669 );
not ( w7197 , w7196 );
and ( w7198 , w7197 , w7038 );
and ( w7199 , w7198 , w7345 );
and ( w7200 , w7199 , g13 );
not ( w7201 , w7200 );
and ( w7202 , w7119 , w7201 );
and ( w7203 , w7202 , g6 );
nor ( w7204 , w7203 , g11 );
and ( w7205 , w7204 , w7345 );
nor ( w7206 , w7205 , w7021 );
and ( w7207 , w7206 , g2 );
and ( w7208 , w7207 , g6 );
not ( w7209 , w7208 );
and ( w7210 , w7209 , g6 );
nor ( w7211 , w7210 , w2669 );
not ( w7212 , w7211 );
and ( w7213 , w7212 , w7038 );
and ( w7214 , w7213 , w7345 );
nor ( w7215 , w7214 , w7021 );
not ( w7216 , w7043 );
and ( w7217 , w7215 , w7216 );
and ( w7218 , w7217 , g2 );
not ( w7219 , w7218 );
and ( w7220 , w7219 , w7113 );
nor ( w7221 , w7220 , w7021 );
and ( w7222 , w7221 , w8382 );
and ( w7223 , w7222 , g14 );
not ( w7224 , w7223 );
and ( w7225 , w7224 , w7038 );
and ( w7226 , w7225 , w7345 );
not ( w7227 , w7226 );
and ( w7228 , w7227 , g17 );
not ( w7229 , w7228 );
and ( w7230 , w7229 , w7039 );
nor ( w7231 , w7230 , g11 );
not ( w7232 , w7231 );
and ( w7233 , w7232 , w7039 );
and ( w7234 , w7233 , g6 );
nor ( w7235 , w7234 , w2669 );
not ( w7236 , w7235 );
and ( w7237 , w7236 , w7038 );
and ( w7238 , w7237 , w7345 );
not ( w7239 , w7238 );
and ( w7240 , w7239 , g2 );
not ( w7241 , w7240 );
and ( w7242 , w7241 , w7113 );
nor ( w7243 , w7069 , w7242 );
and ( w7244 , w7243 , w7044 );
not ( w7245 , w7244 );
and ( w7246 , w7245 , g13 );
not ( w7247 , w7246 );
and ( w7248 , w7247 , g6 );
and ( w7249 , w7248 , w7783 );
and ( w7250 , w7249 , w8382 );
and ( w7251 , w7250 , g14 );
not ( w7252 , w7251 );
and ( w7253 , w7252 , w7039 );
and ( w7254 , w7044 , w8382 );
and ( w7255 , w7254 , g14 );
and ( w7256 , w7255 , g2 );
not ( w7257 , w7256 );
and ( w7258 , w7253 , w7257 );
not ( w7259 , w7258 );
and ( w7260 , w7259 , g3 );
nor ( w7261 , w7260 , w7020 );
and ( w7262 , w7261 , w7039 );
not ( w7263 , w7262 );
and ( w7264 , w7263 , g6 );
not ( w7265 , w7264 );
and ( w7266 , w7265 , w7038 );
and ( w7267 , w7143 , g12 );
and ( w7268 , w7267 , w8382 );
and ( w7269 , w7268 , g14 );
and ( w7270 , w7269 , w8860 );
and ( w7271 , w7270 , w8730 );
nor ( w7272 , w7271 , w7020 );
and ( w7273 , w7272 , w7038 );
not ( w7274 , w7273 );
and ( w7275 , w7274 , g2 );
not ( w7276 , w7275 );
and ( w7277 , w7276 , w7039 );
nor ( w7278 , w7277 , g6 );
not ( w7279 , w7278 );
and ( w7280 , w7279 , w7038 );
and ( w7281 , w7280 , w7345 );
nor ( w7282 , w7281 , g11 );
nor ( w7283 , w7282 , w7020 );
not ( w7284 , w7283 );
and ( w7285 , w7284 , g17 );
and ( w7286 , w7285 , g3 );
not ( w7287 , w7286 );
and ( w7288 , w7287 , w7039 );
and ( w7289 , w7266 , w7288 );
nor ( w7290 , w7289 , g11 );
nor ( w7291 , w7290 , w7020 );
not ( w7292 , w7291 );
and ( w7293 , w7292 , g17 );
and ( w7294 , w7293 , w4849 );
not ( w7295 , w7294 );
and ( w7296 , w7295 , w7038 );
and ( w7297 , w7296 , w7039 );
and ( w7298 , w7297 , g16 );
nor ( w7299 , w7298 , w7242 );
and ( w7300 , w7299 , w7044 );
not ( w7301 , w7300 );
and ( w7302 , w7301 , g13 );
nor ( w7303 , w7057 , w7302 );
nor ( w7304 , w7303 , w7020 );
not ( w7305 , w7304 );
and ( w7306 , w7305 , g2 );
not ( w7307 , w7306 );
and ( w7308 , w7307 , w7038 );
not ( w7309 , w7308 );
and ( w7310 , w7309 , g2 );
and ( w7311 , w7310 , g6 );
not ( w7312 , w7311 );
and ( w7313 , w7312 , w7038 );
nor ( w7314 , w7313 , g16 );
and ( w7315 , w7314 , g2 );
not ( w7316 , w7315 );
and ( w7317 , w7316 , w7039 );
not ( w7318 , w7317 );
and ( w7319 , w7318 , g11 );
not ( w7320 , w7319 );
and ( w7321 , w7320 , w7039 );
and ( w7322 , w7039 , w8819 );
nor ( w7323 , w7322 , w7302 );
and ( w7324 , w7323 , w7783 );
nor ( w7325 , w7324 , w7020 );
nor ( w7326 , w7325 , g11 );
not ( w7327 , w7326 );
and ( w7328 , w7039 , w7327 );
not ( w7329 , w7328 );
and ( w7330 , w7329 , g6 );
not ( w7331 , w7330 );
and ( w7332 , w7331 , w7038 );
and ( w7333 , w7332 , w7345 );
and ( w7334 , w7044 , w8845 );
and ( w7335 , w7334 , g9 );
nor ( w7336 , w7335 , w7020 );
not ( w7337 , w7336 );
and ( w7338 , w7337 , g1 );
not ( w7339 , w7338 );
and ( w7340 , w7339 , w7038 );
nor ( w7341 , w7340 , g13 );
and ( w7342 , w7341 , w7040 );
not ( w7343 , w7342 );
and ( w7344 , w7343 , w7038 );
not ( w7345 , w7020 );
and ( w7346 , w7344 , w7345 );
nor ( w7347 , w7346 , g6 );
and ( w7348 , w7347 , g2 );
and ( w7349 , w7348 , w8828 );
and ( w7350 , w7349 , g9 );
nor ( w7351 , w7350 , w7020 );
not ( w7352 , w7351 );
and ( w7353 , w7352 , w400 );
not ( w7354 , w7353 );
and ( w7355 , w7039 , w7354 );
not ( w7356 , w7355 );
and ( w7357 , w7356 , g11 );
nor ( w7358 , w7357 , w7323 );
not ( w7359 , w7358 );
and ( w7360 , w7359 , g2 );
and ( w7361 , w7058 , w8845 );
not ( w7362 , w7113 );
and ( w7363 , w7361 , w7362 );
not ( w7364 , w7042 );
and ( w7365 , w7364 , w7363 );
not ( w7366 , w7365 );
and ( w7367 , w7039 , w7366 );
not ( w7368 , w7367 );
and ( w7369 , w7368 , g11 );
not ( w7370 , w7369 );
and ( w7371 , w7370 , w7039 );
and ( w7372 , w7371 , w8819 );
nor ( w7373 , w7372 , w7113 );
and ( w7374 , w7373 , w8828 );
not ( w7375 , w7374 );
and ( w7376 , w7375 , w7038 );
and ( w7377 , w7376 , w7039 );
not ( w7378 , w7360 );
and ( w7379 , w7378 , w7377 );
nor ( w7380 , w7379 , g6 );
not ( w7381 , w7380 );
and ( w7382 , w7333 , w7381 );
and ( w7383 , w7321 , w7382 );
and ( w7384 , w7383 , w8819 );
nor ( w7385 , w7384 , w7302 );
and ( w7386 , w7385 , w8828 );
nor ( w7387 , w7386 , w7020 );
and ( w7388 , w7387 , w7038 );
not ( w7389 , w7388 );
and ( w7390 , w7389 , g2 );
not ( w7391 , w7390 );
and ( w7392 , w7391 , w7038 );
and ( t_10 , w7392 , w7383 );
and ( w7393 , g6 , g11 );
and ( w7394 , w7393 , g16 );
nor ( w7395 , w7394 , g13 );
and ( w7396 , w8382 , g14 );
and ( w7397 , w7396 , w8730 );
and ( w7398 , w7397 , g6 );
and ( w7399 , w7398 , w7783 );
not ( w7400 , w7399 );
and ( w7401 , w7400 , g16 );
nor ( w7402 , w1651 , g6 );
and ( w7403 , w7402 , w8828 );
and ( w7404 , w7403 , w8837 );
and ( w7405 , w7404 , g13 );
nor ( w7406 , w7405 , g16 );
nor ( w7407 , w7401 , w7406 );
and ( w7408 , w7407 , w8837 );
not ( w7409 , w7408 );
and ( w7410 , w7409 , g13 );
nor ( w7411 , w7410 , g2 );
and ( w7412 , w7411 , g6 );
nor ( w7413 , w2669 , g16 );
and ( w7414 , w7413 , g13 );
and ( w7415 , w7414 , w8845 );
nor ( w7416 , w7412 , w7415 );
not ( w7417 , w7416 );
and ( w7418 , w7417 , g9 );
and ( w7419 , w7418 , g1 );
and ( w7420 , w7419 , g3 );
not ( w7421 , w7420 );
and ( w7422 , w7421 , g17 );
and ( w7423 , w7422 , g1 );
and ( w7424 , w7423 , g3 );
and ( w7425 , w7424 , g9 );
nor ( w7426 , w7425 , g2 );
not ( w7427 , w7426 );
and ( w7428 , w7427 , g13 );
not ( w7429 , w7428 );
and ( w7430 , w7429 , g1 );
and ( w7431 , w7430 , g3 );
and ( w7432 , w7431 , g9 );
not ( w7433 , w7432 );
and ( w7434 , w7433 , g17 );
and ( w7435 , w7434 , g1 );
and ( w7436 , w7435 , g3 );
and ( w7437 , w7436 , g9 );
nor ( w7438 , w7437 , g2 );
not ( w7439 , w7395 );
and ( w7440 , w7439 , w7438 );
and ( w7441 , w7440 , g1 );
and ( w7442 , w7441 , g3 );
and ( w7443 , w7442 , g9 );
not ( w7444 , w7443 );
and ( w7445 , w7444 , g17 );
and ( w7446 , w7445 , g1 );
and ( w7447 , w7446 , g3 );
and ( w7448 , w7447 , g9 );
not ( w7449 , w1588 );
and ( w7450 , w7449 , g9 );
and ( w7451 , w7450 , w4849 );
and ( w7452 , w8260 , g13 );
and ( w7453 , w7452 , g9 );
not ( w7454 , w7453 );
and ( w7455 , w7454 , g1 );
not ( w7456 , w7455 );
and ( w7457 , w7456 , g13 );
and ( w7458 , w104 , g16 );
and ( w7459 , w7458 , g8 );
nor ( w7460 , w7459 , g13 );
nor ( w7461 , w7460 , g2 );
not ( w7462 , w7457 );
and ( w7463 , w7462 , w7461 );
and ( w7464 , w7463 , w8845 );
not ( w7465 , w7464 );
and ( w7466 , w7465 , g9 );
not ( w7467 , w7466 );
and ( w7468 , w7467 , g1 );
and ( w7469 , w7468 , w7783 );
nor ( w7470 , g6 , w7469 );
not ( w7471 , w7470 );
and ( w7472 , w7471 , g9 );
not ( w7473 , w7472 );
and ( w7474 , w7473 , g9 );
and ( w7475 , g16 , w8819 );
and ( w7476 , w7451 , g17 );
nor ( w7477 , w7475 , w7476 );
and ( w7478 , w7477 , g9 );
not ( w7479 , w7478 );
and ( w7480 , w7479 , g6 );
nor ( w7481 , w4833 , g2 );
not ( w7482 , w7481 );
and ( w7483 , w7482 , g9 );
not ( w7484 , w7483 );
and ( w7485 , w7484 , g9 );
nor ( w7486 , w7485 , g6 );
nor ( w7487 , w7486 , g6 );
and ( w7488 , w7487 , g8 );
and ( w7489 , w7488 , w7973 );
nor ( w7490 , w7489 , g13 );
nor ( w7491 , w7490 , g2 );
and ( w7492 , w7491 , w104 );
not ( w7493 , w7492 );
and ( w7494 , w7493 , g11 );
nor ( w7495 , g16 , w7494 );
not ( w7496 , w7495 );
and ( w7497 , w7496 , g9 );
and ( w7498 , w7497 , w8819 );
and ( w7499 , g17 , g9 );
and ( w7500 , w7499 , w4849 );
not ( w7501 , w7500 );
and ( w7502 , w7501 , g9 );
and ( w7503 , w7502 , g13 );
not ( w7504 , w7503 );
and ( w7505 , w7504 , g1 );
not ( w7506 , w7498 );
and ( w7507 , w7506 , w7505 );
and ( w7508 , w7507 , w8845 );
not ( w7509 , w7508 );
and ( w7510 , w7509 , g11 );
nor ( w7511 , w7510 , g2 );
nor ( w7512 , w7480 , w7511 );
not ( w7513 , w7512 );
and ( w7514 , w7513 , g1 );
not ( w7515 , w7514 );
and ( w7516 , w7515 , g11 );
nor ( w7517 , w7516 , g2 );
not ( w7518 , w7474 );
and ( w7519 , w7518 , w7517 );
and ( w7520 , w7519 , g1 );
nor ( w7521 , w3323 , g6 );
and ( w7522 , w1414 , g17 );
not ( w7523 , w7522 );
and ( w7524 , w1431 , w7523 );
not ( w7525 , w7524 );
and ( w7526 , w7525 , g6 );
and ( w7527 , w7526 , g13 );
not ( w7528 , w7527 );
and ( w7529 , w7528 , g9 );
not ( w7530 , w7529 );
and ( w7531 , w7530 , g14 );
and ( w7532 , w7531 , w8168 );
nor ( w7533 , w7532 , g1 );
not ( w7534 , w7521 );
and ( w7535 , w7534 , w7533 );
and ( w7536 , w7535 , g9 );
nor ( w7537 , w3655 , g5 );
nor ( w7538 , w7537 , g9 );
and ( w7539 , w7538 , w8792 );
and ( w7540 , w7539 , g2 );
not ( w7541 , w7540 );
and ( w7542 , w7541 , g2 );
nor ( w7543 , w7542 , g4 );
and ( w7544 , w7543 , w8735 );
and ( w7545 , w7544 , w8792 );
nor ( w7546 , w3736 , g3 );
and ( w7547 , w467 , w7546 );
and ( w7548 , w7547 , w8765 );
and ( w7549 , w7548 , w8792 );
not ( w7550 , w7549 );
and ( w7551 , w7550 , g2 );
not ( w7552 , w7551 );
and ( w7553 , w7552 , g4 );
and ( w7554 , w7553 , w8845 );
and ( w7555 , w7554 , w8735 );
and ( w7556 , w7555 , w408 );
nor ( w7557 , w7556 , g1 );
not ( w7558 , w7545 );
and ( w7559 , w7558 , w7557 );
nor ( w7560 , w7559 , g3 );
and ( w7561 , w7560 , w8845 );
nor ( w7562 , w7561 , g3 );
and ( w7563 , w7562 , w8765 );
nor ( w7564 , w7563 , g1 );
nor ( w7565 , w7564 , g1 );
nor ( w7566 , g3 , w7565 );
and ( w7567 , w3656 , w8767 );
and ( w7568 , w7567 , g12 );
and ( w7569 , w7568 , w8742 );
nor ( w7570 , w7566 , w7569 );
not ( w7571 , w7570 );
and ( w7572 , w7571 , g13 );
not ( w7573 , w7572 );
and ( w7574 , w7573 , g6 );
nor ( w7575 , w7574 , w42 );
nor ( w7576 , w7575 , g9 );
and ( w7577 , w7576 , w7783 );
not ( w7578 , w7577 );
and ( w7579 , w7578 , g14 );
and ( w7580 , w7579 , w8168 );
and ( w7581 , w290 , g6 );
nor ( w7582 , w7581 , w5038 );
not ( w7583 , w7582 );
and ( w7584 , w7583 , g6 );
nor ( w7585 , w7584 , w471 );
nor ( w7586 , w7585 , g9 );
and ( w7587 , w7586 , w8792 );
and ( w7588 , w526 , w7587 );
and ( w7589 , w8765 , g7 );
nor ( w7590 , w7589 , w59 );
and ( w7591 , w7590 , w8769 );
nor ( w7592 , w7591 , g6 );
and ( w7593 , w2001 , g5 );
and ( w7594 , w7593 , w8845 );
not ( w7595 , w7594 );
and ( w7596 , w7595 , g5 );
nor ( w7597 , w7596 , g4 );
and ( w7598 , w7597 , w8845 );
and ( w7599 , w7598 , w8792 );
and ( w7600 , w7592 , w7599 );
nor ( w7601 , w6890 , w7600 );
nor ( w7602 , w7601 , w3526 );
nor ( w7603 , w7602 , g12 );
and ( w7604 , w4879 , g3 );
and ( w7605 , w7604 , w8792 );
not ( w7606 , w7603 );
and ( w7607 , w7606 , w7605 );
and ( w7608 , w7607 , w8845 );
nor ( w7609 , w7608 , w381 );
not ( w7610 , w7609 );
and ( w7611 , w7610 , g3 );
nor ( w7612 , w7611 , g16 );
nor ( w7613 , w7612 , g1 );
not ( w7614 , w7613 );
and ( w7615 , w7614 , g11 );
not ( w7616 , w7588 );
and ( w7617 , w7616 , w7615 );
not ( w7618 , w7617 );
and ( w7619 , w7618 , g3 );
and ( w7620 , w7619 , w8792 );
and ( w7621 , w7620 , w7783 );
and ( w7622 , w5819 , w7621 );
not ( w7623 , w3320 );
and ( w7624 , w7623 , g9 );
and ( w7625 , w7624 , w7783 );
nor ( w7626 , w7622 , w7625 );
not ( w7627 , w7626 );
and ( w7628 , w7627 , g3 );
and ( w7629 , w1720 , w8765 );
not ( w7630 , w7629 );
and ( w7631 , w7630 , w40 );
nor ( w7632 , w7631 , g3 );
nor ( w7633 , w7632 , g2 );
and ( w7634 , w7633 , w8792 );
and ( w7635 , w7634 , w8845 );
not ( w7636 , w7635 );
and ( w7637 , w7636 , g16 );
not ( w7638 , w7637 );
and ( w7639 , w7638 , w104 );
and ( w7640 , w7639 , w7997 );
and ( w7641 , w7640 , w8792 );
nor ( w7642 , w7641 , g11 );
not ( w7643 , w7642 );
and ( w7644 , w7643 , g13 );
not ( w7645 , w7644 );
and ( w7646 , g10 , w7645 );
not ( w7647 , w7646 );
and ( w7648 , w7647 , g9 );
and ( w7649 , w8792 , w361 );
nor ( w7650 , w7649 , g3 );
not ( w7651 , w7650 );
and ( w7652 , w7651 , g4 );
and ( w7653 , w7652 , w7783 );
and ( w7654 , w7653 , w8845 );
and ( w7655 , w7654 , w4833 );
nor ( w7656 , w7655 , w4977 );
not ( w7657 , w7656 );
and ( w7658 , w7657 , w408 );
and ( w7659 , w7658 , w8730 );
not ( w7660 , w7659 );
and ( w7661 , w7660 , g14 );
and ( w7662 , w7661 , w8168 );
nor ( w7663 , w381 , g12 );
and ( w7664 , w7663 , g4 );
and ( w7665 , w7664 , w8769 );
and ( w7666 , w7665 , w8742 );
not ( w7667 , w7666 );
and ( w7668 , w7667 , w40 );
nor ( w7669 , w7668 , w4954 );
nor ( w7670 , w7669 , g2 );
and ( w7671 , w7670 , w8792 );
not ( w7672 , w7662 );
and ( w7673 , w7672 , w7671 );
and ( w7674 , w7673 , w408 );
and ( w7675 , w7674 , w8845 );
not ( w7676 , w7675 );
and ( w7677 , w7676 , g16 );
not ( w7678 , w7677 );
and ( w7679 , w7678 , w104 );
not ( w7680 , w7679 );
and ( w7681 , w7680 , g13 );
not ( w7682 , w7681 );
and ( w7683 , w7682 , w104 );
and ( w7684 , w7683 , w8792 );
nor ( w7685 , w7684 , g11 );
not ( w7686 , w7648 );
and ( w7687 , w7686 , w7685 );
and ( w7688 , w7687 , g16 );
not ( w7689 , w7688 );
and ( w7690 , w7689 , w104 );
not ( w7691 , w7690 );
and ( w7692 , w7691 , g13 );
nor ( w7693 , w7692 , g2 );
and ( w7694 , w7693 , w8845 );
and ( w7695 , w7694 , w8792 );
nor ( w7696 , w2022 , w7695 );
nor ( w7697 , w2191 , g4 );
and ( w7698 , w7697 , w8769 );
nor ( w7699 , w7698 , g3 );
nor ( w7700 , w7699 , g7 );
and ( w7701 , w7700 , g8 );
and ( w7702 , w8765 , w7701 );
nor ( w7703 , w7696 , w7702 );
and ( w7704 , w7703 , w8735 );
nor ( w7705 , w7628 , w7704 );
and ( w7706 , w7705 , w8819 );
nor ( w7707 , w7706 , w7696 );
not ( w7708 , w7580 );
and ( w7709 , w7708 , w7707 );
not ( w7710 , w7709 );
and ( w7711 , w7710 , g16 );
not ( w7712 , w7711 );
and ( w7713 , w7712 , w7707 );
not ( w7714 , w7713 );
and ( w7715 , w7714 , g11 );
and ( w7716 , w7783 , w2619 );
nor ( w7717 , w7716 , w104 );
and ( w7718 , w7717 , w7783 );
and ( w7719 , w408 , g3 );
and ( w7720 , w7719 , w1489 );
nor ( w7721 , w7720 , w104 );
not ( w7722 , w7721 );
and ( w7723 , w7722 , g3 );
nor ( w7724 , w7718 , w7723 );
not ( w7725 , w104 );
and ( w7726 , w7724 , w7725 );
nor ( w7727 , w7726 , w7696 );
and ( w7728 , w7727 , g3 );
nor ( w7729 , w7704 , g13 );
nor ( w7730 , w7729 , g2 );
nor ( w7731 , w7728 , w7730 );
nor ( w7732 , w6323 , g10 );
and ( w7733 , w7732 , w8767 );
nor ( w7734 , w7733 , g6 );
and ( w7735 , w7734 , g9 );
nor ( w7736 , g6 , w7735 );
not ( w7737 , w7736 );
and ( w7738 , w7737 , g9 );
nor ( w7739 , w5377 , g4 );
and ( w7740 , w7739 , w8769 );
and ( w7741 , w7740 , w8742 );
and ( w7742 , w7741 , g8 );
not ( w7743 , w7742 );
and ( w7744 , w7743 , w33 );
not ( w7745 , w7744 );
and ( w7746 , w7745 , g10 );
nor ( w7747 , w7746 , g6 );
and ( w7748 , w7747 , w8735 );
nor ( w7749 , g6 , w7748 );
nor ( w7750 , w7749 , g9 );
and ( w7751 , w7750 , w8735 );
nor ( w7752 , w7738 , w7751 );
nor ( w7753 , w41 , g9 );
nor ( w7754 , w7753 , g3 );
and ( w7755 , w7754 , w7783 );
not ( w7756 , w7752 );
and ( w7757 , w7756 , w7755 );
nor ( w7758 , w467 , w2687 );
nor ( w7759 , w7758 , g9 );
and ( w7760 , w7759 , g3 );
and ( w7761 , w7760 , w8845 );
nor ( w7762 , w7761 , w7735 );
and ( w7763 , w8845 , w7762 );
nor ( w7764 , w5929 , g9 );
and ( w7765 , w2026 , w8769 );
and ( w7766 , w7765 , w8765 );
and ( w7767 , w7766 , w1984 );
nor ( w7768 , w7767 , g7 );
and ( w7769 , w7768 , w8860 );
and ( w7770 , w7769 , w8769 );
not ( w7771 , w7770 );
and ( w7772 , w7764 , w7771 );
and ( w7773 , w7772 , g6 );
and ( w7774 , w7773 , w8792 );
nor ( w7775 , g9 , w7774 );
not ( w7776 , w7775 );
and ( w7777 , w7776 , w1489 );
nor ( w7778 , w3371 , w7761 );
not ( w7779 , w7777 );
and ( w7780 , w7779 , w7778 );
not ( w7781 , w7780 );
and ( w7782 , w7781 , g3 );
not ( w7783 , g2 );
and ( w7784 , w7782 , w7783 );
not ( w7785 , w7763 );
and ( w7786 , w7785 , w7784 );
nor ( w7787 , w7757 , w7786 );
nor ( w7788 , w7695 , g16 );
and ( w7789 , w7788 , w8819 );
nor ( w7790 , w7789 , g2 );
nor ( w7791 , w2022 , w7790 );
nor ( w7792 , w7787 , w7791 );
nor ( w7793 , w7792 , g16 );
nor ( w7794 , w7793 , g2 );
not ( w7795 , w7731 );
and ( w7796 , w7795 , w7794 );
nor ( w7797 , w7796 , g13 );
nor ( w7798 , w7502 , g2 );
not ( w7799 , w7798 );
and ( w7800 , w7799 , g16 );
nor ( w7801 , w7800 , w7406 );
and ( w7802 , w7801 , g1 );
and ( w7803 , w7696 , g13 );
and ( w7804 , w7803 , w8837 );
nor ( w7805 , w7804 , g2 );
nor ( w7806 , w7802 , w7805 );
nor ( w7807 , w7797 , w7806 );
nor ( w7808 , w7807 , g11 );
nor ( w7809 , w7808 , g2 );
not ( w7810 , w7715 );
and ( w7811 , w7810 , w7809 );
nor ( w7812 , w7536 , w7811 );
nor ( w7813 , w7812 , g2 );
and ( w7814 , w7813 , w7707 );
not ( w7815 , w7814 );
and ( w7816 , w7815 , g11 );
not ( w7817 , w7816 );
and ( w7818 , w7817 , w7809 );
nor ( w7819 , w7520 , w7818 );
and ( w7820 , w7819 , g11 );
not ( w7821 , w7820 );
and ( w7822 , w7821 , w7809 );
not ( w7823 , w7448 );
and ( w7824 , w7823 , w7822 );
and ( w7825 , w7040 , g11 );
nor ( w7826 , w7825 , g13 );
not ( w7827 , w7826 );
and ( w7828 , w7827 , g9 );
and ( w7829 , w7828 , w4912 );
and ( w7830 , g2 , w8765 );
nor ( w7831 , w7830 , w7824 );
nor ( w7832 , w7831 , g9 );
and ( w7833 , w7832 , g11 );
not ( w7834 , w7450 );
and ( w7835 , w7834 , g1 );
and ( w7836 , w7499 , w8730 );
and ( w7837 , g9 , g10 );
nor ( w7838 , w7837 , w7569 );
and ( w7839 , w7838 , w408 );
and ( w7840 , w7839 , g11 );
not ( w7841 , w7840 );
and ( w7842 , w7841 , g13 );
not ( w7843 , w7842 );
and ( w7844 , w7843 , g2 );
nor ( w7845 , w7844 , w7824 );
not ( w7846 , w7836 );
and ( w7847 , w7846 , w7845 );
not ( w7848 , w7847 );
and ( w7849 , w7848 , w1473 );
not ( w7850 , w1430 );
and ( w7851 , w7850 , w7845 );
not ( w7852 , w7851 );
and ( w7853 , w7852 , w381 );
and ( w7854 , w7853 , g16 );
nor ( w7855 , w5802 , g1 );
nor ( w7856 , g2 , w7824 );
and ( w7857 , w7855 , w8274 );
and ( w7858 , w7857 , g9 );
nor ( w7859 , w5118 , w7824 );
nor ( w7860 , w3947 , w7859 );
and ( w7861 , w7860 , g3 );
and ( w7862 , w7861 , w8833 );
nor ( w7863 , w7862 , g15 );
and ( w7864 , w1536 , g12 );
and ( w7865 , w7864 , w27 );
nor ( w7866 , w4954 , w7865 );
nor ( w7867 , w7866 , g4 );
nor ( w7868 , w1846 , w7824 );
not ( w7869 , w7867 );
and ( w7870 , w7869 , w7868 );
nor ( w7871 , w7870 , g10 );
and ( w7872 , w7871 , w8792 );
and ( w7873 , w7872 , g2 );
and ( w7874 , w7873 , g11 );
nor ( w7875 , w2896 , g18 );
and ( w7876 , w7875 , g9 );
and ( w7877 , w7876 , w8860 );
and ( w7878 , w7877 , g17 );
and ( w7879 , w7878 , g12 );
and ( w7880 , w7879 , g14 );
and ( w7881 , w7880 , w8730 );
and ( w7882 , w7881 , g16 );
nor ( w7883 , w7882 , w7405 );
not ( w7884 , w7883 );
and ( w7885 , w7884 , g9 );
not ( w7886 , w7885 );
and ( w7887 , w7886 , w7831 );
not ( w7888 , w7887 );
and ( w7889 , w7888 , w4849 );
not ( w7890 , w1981 );
and ( w7891 , w7890 , g2 );
and ( w7892 , w7891 , w8765 );
and ( w7893 , w7892 , w8735 );
nor ( w7894 , w7893 , w7824 );
not ( w7895 , w7889 );
and ( w7896 , w7895 , w7894 );
not ( w7897 , w7896 );
and ( w7898 , w7897 , g1 );
and ( w7899 , w7898 , w8837 );
not ( w7900 , w7899 );
and ( w7901 , w7900 , g13 );
not ( w7902 , w7901 );
and ( w7903 , w7902 , g2 );
and ( w7904 , w7903 , g1 );
nor ( w7905 , w241 , w7824 );
not ( w7906 , w7904 );
and ( w7907 , w7906 , w7905 );
nor ( w7908 , w7907 , g11 );
and ( w7909 , w7908 , w400 );
not ( w7910 , w7909 );
and ( w7911 , w7910 , g13 );
not ( w7912 , w7911 );
and ( w7913 , w7912 , g2 );
nor ( w7914 , w7913 , w7824 );
not ( w7915 , w7874 );
and ( w7916 , w7915 , w7914 );
nor ( w7917 , w7916 , g6 );
and ( w7918 , w7917 , g2 );
nor ( w7919 , w7918 , w7824 );
nor ( w7920 , w7863 , w7919 );
not ( w7921 , w7865 );
and ( w7922 , w7921 , w7868 );
nor ( w7923 , w7922 , g3 );
and ( w7924 , w7923 , w8792 );
and ( w7925 , w7924 , g2 );
and ( w7926 , w7925 , g11 );
not ( w7927 , w7926 );
and ( w7928 , w7927 , w7914 );
nor ( w7929 , w7928 , g6 );
and ( w7930 , w7929 , g2 );
nor ( w7931 , w7930 , w7824 );
not ( w7932 , w7920 );
and ( w7933 , w7932 , w7931 );
not ( w7934 , w381 );
and ( w7935 , w7933 , w7934 );
nor ( w7936 , w7935 , g10 );
and ( w7937 , w7936 , w8765 );
and ( w7938 , w7937 , w8792 );
and ( w7939 , w7938 , g11 );
not ( w7940 , w7939 );
and ( w7941 , w7940 , w7914 );
nor ( w7942 , w7941 , g6 );
and ( w7943 , w7942 , g2 );
nor ( w7944 , w7943 , w7824 );
not ( w7945 , w7944 );
and ( w7946 , w1408 , w7945 );
and ( w7947 , w7860 , g10 );
and ( w7948 , w7947 , g3 );
not ( w7949 , w7948 );
and ( w7950 , w7949 , w7931 );
nor ( w7951 , w7950 , w213 );
and ( w7952 , w7951 , g10 );
and ( w7953 , w7952 , w8792 );
and ( w7954 , w7953 , g11 );
not ( w7955 , w7954 );
and ( w7956 , w7955 , w7914 );
nor ( w7957 , w7956 , g6 );
and ( w7958 , w7957 , g2 );
nor ( w7959 , w7958 , w7824 );
not ( w7960 , w7946 );
and ( w7961 , w7960 , w7959 );
nor ( w7962 , w7961 , g9 );
and ( w7963 , w7962 , w8792 );
and ( w7964 , w7963 , g11 );
not ( w7965 , w7964 );
and ( w7966 , w7965 , w7914 );
not ( w7967 , w7858 );
and ( w7968 , w7967 , w7966 );
and ( w7969 , w213 , g9 );
and ( w7970 , w7969 , g8 );
and ( w7971 , w7970 , w8730 );
nor ( w7972 , w7968 , w7971 );
not ( w7973 , g17 );
and ( w7974 , w7972 , w7973 );
not ( w7975 , w76 );
and ( w7976 , w7975 , w213 );
nor ( w7977 , w7976 , w7856 );
and ( w7978 , w7977 , g9 );
and ( w7979 , w1350 , w8730 );
and ( w7980 , w7979 , w381 );
not ( w7981 , w7868 );
and ( w7982 , w7981 , g4 );
and ( w7983 , w1264 , w8769 );
nor ( w7984 , w7983 , w7831 );
and ( w7985 , w7984 , g3 );
and ( w7986 , w7985 , w8765 );
and ( w7987 , w7986 , w2687 );
nor ( w7988 , w7982 , w7987 );
not ( w7989 , w7988 );
and ( w7990 , w7989 , g3 );
not ( w7991 , w7990 );
and ( w7992 , w7991 , w7931 );
nor ( w7993 , w7992 , g15 );
nor ( w7994 , w7993 , g15 );
and ( w7995 , w7994 , w8382 );
nor ( w7996 , w7995 , w7919 );
not ( w7997 , w213 );
and ( w7998 , w7996 , w7997 );
and ( w7999 , w7998 , w8730 );
and ( w8000 , w7999 , g17 );
and ( w8001 , w8000 , w8792 );
and ( w8002 , w8001 , g11 );
not ( w8003 , w8002 );
and ( w8004 , w8003 , w7914 );
nor ( w8005 , w8004 , g6 );
and ( w8006 , w8005 , g2 );
nor ( w8007 , w8006 , w7824 );
not ( w8008 , w7980 );
and ( w8009 , w8008 , w8007 );
nor ( w8010 , w8009 , g10 );
and ( w8011 , w8010 , g17 );
and ( w8012 , w8011 , w8792 );
and ( w8013 , w8012 , g11 );
not ( w8014 , w8013 );
and ( w8015 , w8014 , w7914 );
nor ( w8016 , w8015 , g6 );
and ( w8017 , w8016 , g2 );
nor ( w8018 , w8017 , w7824 );
and ( w8019 , w8018 , w7959 );
not ( w8020 , w8019 );
and ( w8021 , w8020 , g17 );
and ( w8022 , w8021 , w8792 );
not ( w8023 , w8022 );
and ( w8024 , w8023 , w7914 );
not ( w8025 , w7978 );
and ( w8026 , w8025 , w8024 );
not ( w8027 , w8026 );
and ( w8028 , w8027 , g17 );
and ( w8029 , w8028 , w8792 );
and ( w8030 , w8029 , g11 );
not ( w8031 , w8030 );
and ( w8032 , w8031 , w7914 );
nor ( w8033 , w8032 , g6 );
and ( w8034 , w8033 , g2 );
nor ( w8035 , w8034 , w7824 );
not ( w8036 , w7974 );
and ( w8037 , w8036 , w8035 );
nor ( w8038 , w8037 , g16 );
and ( w8039 , w8038 , w8792 );
and ( w8040 , w8039 , g11 );
not ( w8041 , w8040 );
and ( w8042 , w8041 , w7914 );
nor ( w8043 , w8042 , g6 );
not ( w8044 , w8043 );
and ( w8045 , w8044 , g13 );
not ( w8046 , w8045 );
and ( w8047 , w8046 , g2 );
nor ( w8048 , w8047 , w7824 );
not ( w8049 , w7854 );
and ( w8050 , w8049 , w8048 );
nor ( w8051 , w8050 , g1 );
and ( w8052 , w8051 , g11 );
not ( w8053 , w8052 );
and ( w8054 , w8053 , w7914 );
not ( w8055 , w8054 );
and ( w8056 , w8055 , w400 );
not ( w8057 , w8056 );
and ( w8058 , w8057 , g13 );
not ( w8059 , w8058 );
and ( w8060 , w8059 , g2 );
nor ( w8061 , w8060 , w7824 );
and ( w8062 , w8061 , g13 );
not ( w8063 , w7849 );
and ( w8064 , w8063 , w8062 );
not ( w8065 , w8064 );
and ( w8066 , w8065 , w400 );
not ( w8067 , w8066 );
and ( w8068 , w8067 , g11 );
nor ( w8069 , w1981 , g5 );
and ( w8070 , w8069 , w8742 );
nor ( w8071 , w8070 , g7 );
and ( w8072 , w8071 , w8769 );
not ( w8073 , w8072 );
and ( w8074 , w8073 , g2 );
and ( w8075 , w8074 , w8767 );
nor ( w8076 , w8075 , g8 );
nor ( w8077 , w8076 , g9 );
nor ( w8078 , w1408 , g16 );
nor ( w8079 , w8078 , g9 );
not ( w8080 , w8079 );
and ( w8081 , w8080 , g13 );
not ( w8082 , w8081 );
and ( w8083 , w8082 , w361 );
and ( w8084 , w8083 , w6728 );
not ( w8085 , w8084 );
and ( w8086 , w8085 , g14 );
and ( w8087 , w8086 , w8168 );
not ( w8088 , w8087 );
and ( w8089 , w8088 , g2 );
and ( w8090 , w8089 , g6 );
nor ( w8091 , w8090 , w2022 );
nor ( w8092 , w6716 , g9 );
and ( w8093 , w8092 , g2 );
and ( w8094 , w8093 , w8792 );
and ( w8095 , w8094 , g6 );
and ( w8096 , w8095 , w8079 );
not ( w8097 , w8096 );
and ( w8098 , w8097 , g13 );
nor ( w8099 , w8098 , g3 );
not ( w8100 , w8099 );
and ( w8101 , w8100 , g14 );
and ( w8102 , w8101 , w8168 );
nor ( w8103 , w2441 , w2022 );
not ( w8104 , w4822 );
and ( w8105 , w8104 , w8103 );
nor ( w8106 , w8102 , w8105 );
and ( w8107 , w8106 , w8765 );
and ( w8108 , w8107 , g2 );
nor ( w8109 , w8108 , w2022 );
and ( w8110 , w8109 , w8837 );
not ( w8111 , w8110 );
and ( w8112 , w2441 , w8111 );
nor ( w8113 , w8112 , w2022 );
nor ( w8114 , w8091 , w8113 );
nor ( w8115 , w241 , w7695 );
not ( w8116 , w8114 );
and ( w8117 , w8116 , w8115 );
nor ( w8118 , w8117 , g3 );
and ( w8119 , w8118 , w8765 );
nor ( w8120 , w8119 , g11 );
and ( w8121 , w1588 , w8120 );
nor ( w8122 , w8121 , g3 );
and ( w8123 , w8122 , w8765 );
and ( w8124 , w8077 , w8123 );
and ( w8125 , w8124 , g2 );
nor ( w8126 , w8125 , w7824 );
nor ( w8127 , w8126 , g9 );
and ( w8128 , w8150 , g3 );
not ( w8129 , w8128 );
and ( w8130 , w8129 , w2687 );
nor ( w8131 , w8130 , g4 );
not ( w8132 , w8131 );
and ( w8133 , w8132 , g6 );
and ( w8134 , w8133 , w8792 );
nor ( w8135 , w4449 , w8134 );
and ( w8136 , w8135 , g6 );
and ( w8137 , w1516 , g3 );
not ( w8138 , w8137 );
and ( w8139 , w8138 , w8126 );
nor ( w8140 , w8139 , g1 );
and ( w8141 , g12 , w8767 );
and ( w8142 , w8141 , w8742 );
and ( w8143 , w8142 , w8735 );
and ( w8144 , w8143 , w8860 );
and ( w8145 , w8144 , w8769 );
not ( w8146 , w8145 );
and ( w8147 , w8140 , w8146 );
and ( w8148 , w8147 , g16 );
and ( w8149 , w8148 , w4357 );
not ( w8150 , w4954 );
and ( w8151 , w8150 , w8120 );
nor ( w8152 , w8151 , g9 );
and ( w8153 , w8152 , g16 );
nor ( w8154 , w1366 , w7831 );
and ( w8155 , w8154 , w8828 );
and ( w8156 , w8155 , w8765 );
nor ( w8157 , w8156 , w7824 );
not ( w8158 , w8153 );
and ( w8159 , w8158 , w8157 );
not ( w8160 , w8159 );
and ( w8161 , w8160 , g6 );
and ( w8162 , w8161 , w8730 );
and ( w8163 , w8162 , w8765 );
and ( w8164 , w8163 , g2 );
nor ( w8165 , w8164 , w7824 );
not ( w8166 , w8149 );
and ( w8167 , w8166 , w8165 );
not ( w8168 , w122 );
and ( w8169 , w8167 , w8168 );
and ( w8170 , w8169 , w213 );
nor ( w8171 , w8170 , g9 );
and ( w8172 , w8171 , w8837 );
and ( w8173 , w8172 , g6 );
not ( w8174 , w8173 );
and ( w8175 , w8174 , w8062 );
and ( w8176 , w8175 , g14 );
not ( w8177 , w3370 );
and ( w8178 , w8177 , g6 );
nor ( w8179 , w8178 , g1 );
nor ( w8180 , w8179 , g1 );
not ( w8181 , w8180 );
and ( w8182 , w8181 , g8 );
nor ( w8183 , w8182 , g1 );
and ( w8184 , w8183 , g11 );
and ( w8185 , g10 , g18 );
nor ( w8186 , w8185 , g14 );
not ( w8187 , w8186 );
and ( w8188 , w8187 , g9 );
and ( w8189 , w8188 , g17 );
and ( w8190 , w8189 , g14 );
and ( w8191 , w8190 , w4849 );
nor ( w8192 , w1516 , w8191 );
not ( w8193 , w8192 );
and ( w8194 , w8193 , g2 );
and ( w8195 , w8194 , w8837 );
and ( w8196 , w8195 , g9 );
and ( w8197 , w8196 , g6 );
not ( w8198 , w8197 );
and ( w8199 , w8198 , g13 );
not ( w8200 , w8184 );
and ( w8201 , w8200 , w8199 );
not ( w8202 , w8201 );
and ( w8203 , w8202 , g9 );
not ( w8204 , w8183 );
and ( w8205 , w8204 , g11 );
nor ( w8206 , w6635 , w7824 );
nor ( w8207 , w8205 , w8206 );
and ( w8208 , w8207 , g2 );
not ( w8209 , w8208 );
and ( w8210 , w8209 , w8062 );
nor ( w8211 , w8210 , g9 );
not ( w8212 , w8211 );
and ( w8213 , w8212 , g16 );
not ( w8214 , w8189 );
and ( w8215 , w8214 , g11 );
and ( w8216 , g18 , w8769 );
and ( w8217 , g18 , w8742 );
nor ( w8218 , w8216 , w8217 );
not ( w8219 , w8218 );
and ( w8220 , w8219 , g9 );
and ( w8221 , w8220 , g10 );
nor ( w8222 , w8221 , g14 );
not ( w8223 , w2896 );
and ( w8224 , w8223 , g9 );
and ( w8225 , w8224 , g17 );
not ( w8226 , w8225 );
and ( w8227 , w8226 , g14 );
nor ( w8228 , w8222 , w8227 );
and ( w8229 , w8228 , w8860 );
not ( w8230 , w8229 );
and ( w8231 , w8230 , g12 );
not ( w8232 , w8231 );
and ( w8233 , w8232 , g12 );
and ( w8234 , w8233 , w8274 );
nor ( w8235 , w8234 , g11 );
not ( w8236 , w7824 );
and ( w8237 , w8235 , w8236 );
nor ( w8238 , w8215 , w8237 );
and ( w8239 , w1845 , w4357 );
not ( w8240 , w8239 );
and ( w8241 , w8240 , g10 );
and ( w8242 , w8241 , w8860 );
not ( w8243 , w8242 );
and ( w8244 , w8243 , g3 );
and ( w8245 , w8244 , g9 );
and ( w8246 , w8245 , w4912 );
not ( w8247 , w8246 );
and ( w8248 , w8247 , w7831 );
not ( w8249 , w8248 );
and ( w8250 , w8249 , g2 );
and ( w8251 , w8250 , g6 );
not ( w8252 , w8251 );
and ( w8253 , w8252 , w8062 );
nor ( w8254 , w8253 , g15 );
and ( w8255 , w8254 , g1 );
nor ( w8256 , w1 , w7824 );
not ( w8257 , w8255 );
and ( w8258 , w8257 , w8256 );
and ( w8259 , w8258 , w8828 );
not ( w8260 , w7451 );
and ( w8261 , w8260 , g3 );
not ( w8262 , w8261 );
and ( w8263 , w8262 , w2585 );
not ( w8264 , w8263 );
and ( w8265 , w8264 , w8062 );
not ( w8266 , w8265 );
and ( w8267 , w8266 , g9 );
and ( w8268 , w8267 , g1 );
and ( w8269 , w1473 , w2585 );
not ( w8270 , w8269 );
and ( w8271 , w8270 , g6 );
and ( w8272 , w8271 , w8767 );
nor ( w8273 , w8272 , g1 );
not ( w8274 , w7856 );
and ( w8275 , w8273 , w8274 );
and ( w8276 , w8275 , g9 );
not ( w8277 , w8276 );
and ( w8278 , w8277 , w7831 );
not ( w8279 , w8268 );
and ( w8280 , w8279 , w8278 );
nor ( w8281 , w8280 , w7856 );
not ( w8282 , w8259 );
and ( w8283 , w8282 , w8281 );
not ( w8284 , w8283 );
and ( w8285 , w8284 , g13 );
not ( w8286 , w8285 );
and ( w8287 , w8238 , w8286 );
and ( w8288 , w8287 , w4849 );
and ( w8289 , w8288 , g9 );
not ( w8290 , w8289 );
and ( w8291 , w8290 , w7831 );
not ( w8292 , w8291 );
and ( w8293 , w8292 , g2 );
and ( w8294 , w8293 , g6 );
not ( w8295 , w8294 );
and ( w8296 , w8295 , w8062 );
nor ( w8297 , w8296 , g15 );
and ( w8298 , w8297 , g1 );
not ( w8299 , w8298 );
and ( w8300 , w8299 , w8256 );
and ( w8301 , w8300 , w8828 );
not ( w8302 , w8301 );
and ( w8303 , w8302 , w8281 );
not ( w8304 , w8303 );
and ( w8305 , w8304 , g13 );
nor ( w8306 , w8213 , w8305 );
and ( w8307 , w8306 , w8281 );
and ( w8308 , w8307 , g2 );
nor ( w8309 , w8308 , w7824 );
and ( w8310 , w8309 , g13 );
and ( w8311 , w8310 , w8062 );
and ( w8312 , w6624 , g11 );
and ( w8313 , w8312 , w8792 );
nor ( w8314 , w8313 , w381 );
and ( w8315 , w8314 , g16 );
and ( w8316 , w8315 , g13 );
and ( w8317 , w8311 , w8316 );
nor ( w8318 , w8317 , w8305 );
nor ( w8319 , w8203 , w8318 );
not ( w8320 , w8319 );
and ( w8321 , w8320 , g2 );
and ( w8322 , w8321 , g6 );
not ( w8323 , w8322 );
and ( w8324 , w8323 , w8062 );
and ( w8325 , w8324 , w8316 );
nor ( w8326 , w8325 , w8305 );
not ( w8327 , w8176 );
and ( w8328 , w8327 , w8326 );
nor ( w8329 , w8136 , w8328 );
nor ( w8330 , w8329 , g11 );
and ( w8331 , w8330 , w8765 );
and ( w8332 , w8331 , g6 );
not ( w8333 , w8332 );
and ( w8334 , w8333 , w8062 );
not ( w8335 , w8334 );
and ( w8336 , w8335 , w8326 );
and ( w8337 , w8336 , w8281 );
nor ( w8338 , w8127 , w8337 );
and ( w8339 , w8338 , w8837 );
not ( w8340 , w8339 );
and ( w8341 , w8340 , w8326 );
and ( w8342 , w8341 , w8281 );
not ( w8343 , w8342 );
and ( w8344 , w8343 , g13 );
and ( w8345 , w8360 , w8344 );
nor ( w8346 , w8345 , g1 );
and ( w8347 , w8346 , g6 );
and ( w8348 , w1473 , w8765 );
and ( w8349 , w8348 , w1248 );
and ( w8350 , w8349 , w8735 );
not ( w8351 , w8113 );
and ( w8352 , w8350 , w8351 );
and ( w8353 , w8352 , w1244 );
nor ( w8354 , w8353 , g5 );
and ( w8355 , w8354 , w8765 );
and ( w8356 , w8355 , w8735 );
and ( w8357 , w8356 , w8860 );
and ( w8358 , w8357 , w8742 );
and ( w8359 , w8358 , w8767 );
not ( w8360 , w1431 );
and ( w8361 , w8360 , w8165 );
nor ( w8362 , w8361 , g10 );
and ( w8363 , w8362 , g6 );
and ( w8364 , w8363 , w8792 );
and ( w8365 , w8364 , g2 );
nor ( w8366 , w8365 , w7824 );
and ( w8367 , w8359 , w8366 );
not ( w8368 , w8367 );
and ( w8369 , w8368 , w2585 );
not ( w8370 , w8369 );
and ( w8371 , w8370 , w8115 );
and ( w8372 , w8371 , w8837 );
and ( w8373 , w8372 , g16 );
not ( w8374 , w1347 );
and ( w8375 , w8374 , g11 );
nor ( w8376 , w1517 , w6629 );
not ( w8377 , w8376 );
and ( w8378 , w8377 , g8 );
and ( w8379 , w8378 , w1361 );
and ( w8380 , w8379 , w8382 );
and ( w8381 , w8380 , g3 );
not ( w8382 , g18 );
and ( w8383 , w7971 , w8382 );
and ( w8384 , w8383 , g3 );
not ( w8385 , w8384 );
and ( w8386 , w1353 , w8385 );
and ( w8387 , w8386 , g6 );
nor ( w8388 , w8387 , g11 );
nor ( w8389 , w8388 , g10 );
nor ( w8390 , w8389 , w122 );
nor ( w8391 , w8390 , g1 );
and ( w8392 , w8391 , g2 );
and ( w8393 , w8392 , g6 );
nor ( w8394 , w8393 , w7824 );
not ( w8395 , w8381 );
and ( w8396 , w8395 , w8394 );
nor ( w8397 , w8396 , g10 );
not ( w8398 , w8120 );
and ( w8399 , w8398 , w33 );
nor ( w8400 , w8399 , g9 );
and ( w8401 , w8400 , w8735 );
and ( w8402 , w8401 , g10 );
not ( w8403 , w8402 );
and ( w8404 , w8403 , g6 );
not ( w8405 , w8404 );
and ( w8406 , w8405 , w8115 );
and ( w8407 , w8406 , w213 );
not ( w8408 , w8407 );
and ( w8409 , w8408 , w8326 );
and ( w8410 , w8452 , w8409 );
not ( w8411 , w8410 );
and ( w8412 , w8411 , w8115 );
and ( w8413 , w8412 , w8837 );
and ( w8414 , w8413 , w8828 );
and ( w8415 , w8414 , w213 );
nor ( w8416 , w8415 , g1 );
not ( w8417 , w8416 );
and ( w8418 , w8417 , g14 );
not ( w8419 , w8418 );
and ( w8420 , w8419 , w8326 );
and ( w8421 , w8420 , g2 );
nor ( w8422 , w8421 , w7824 );
and ( w8423 , w8422 , g13 );
not ( w8424 , w8397 );
and ( w8425 , w8424 , w8423 );
not ( w8426 , w8425 );
and ( w8427 , w8426 , w8409 );
and ( w8428 , w8427 , g2 );
and ( w8429 , w8428 , g6 );
not ( w8430 , w8429 );
and ( w8431 , w8430 , w8115 );
and ( w8432 , w8431 , w213 );
nor ( w8433 , w8432 , g1 );
not ( w8434 , w8433 );
and ( w8435 , w8434 , g14 );
not ( w8436 , w8435 );
and ( w8437 , w8436 , w8326 );
and ( w8438 , w8437 , w8281 );
and ( w8439 , w8438 , g2 );
nor ( w8440 , w8439 , w7824 );
and ( w8441 , w8440 , w8115 );
and ( w8442 , w8441 , w8837 );
and ( w8443 , w8442 , w8828 );
and ( w8444 , w8443 , w213 );
not ( w8445 , w8444 );
and ( w8446 , w8445 , w8326 );
not ( w8447 , w8446 );
and ( w8448 , w8447 , g13 );
nor ( w8449 , w8375 , w8448 );
nor ( w8450 , w1517 , w7824 );
nor ( w8451 , g10 , w8450 );
not ( w8452 , w8394 );
and ( w8453 , w8451 , w8452 );
not ( w8454 , w8453 );
and ( w8455 , w8454 , w213 );
nor ( w8456 , w8455 , g1 );
and ( w8457 , w8456 , g2 );
and ( w8458 , w8457 , w8828 );
and ( w8459 , w8458 , g9 );
nor ( w8460 , w5819 , w2585 );
not ( w8461 , w8460 );
and ( w8462 , w8461 , g6 );
and ( w8463 , w8462 , w8765 );
and ( w8464 , w8463 , g6 );
and ( w8465 , w8464 , w8730 );
and ( w8466 , w8465 , w8828 );
and ( w8467 , w8466 , g2 );
nor ( w8468 , w8467 , w7824 );
and ( w8469 , w8468 , w213 );
and ( w8470 , w213 , w8792 );
and ( w8471 , w8470 , g10 );
and ( w8472 , w8471 , w8828 );
nor ( w8473 , w8469 , w8472 );
and ( w8474 , w8473 , g2 );
nor ( w8475 , w8474 , w7824 );
and ( w8476 , w8560 , w8475 );
not ( w8477 , w8476 );
and ( w8478 , w8477 , g6 );
nor ( w8479 , w8478 , g16 );
nor ( w8480 , w8479 , w7831 );
and ( w8481 , w8480 , g11 );
nor ( w8482 , w8481 , w8337 );
nor ( w8483 , w8482 , g9 );
not ( w8484 , w8472 );
and ( w8485 , w8483 , w8484 );
and ( w8486 , w8485 , g6 );
not ( w8487 , w8486 );
and ( w8488 , w8487 , w8062 );
not ( w8489 , w8488 );
and ( w8490 , w8489 , w8326 );
nor ( w8491 , w8459 , w8490 );
not ( w8492 , w8449 );
and ( w8493 , w8492 , w8491 );
not ( w8494 , w8493 );
and ( w8495 , w8494 , g2 );
nor ( w8496 , w8495 , g16 );
and ( w8497 , w8496 , w213 );
and ( w8498 , w8497 , w8597 );
not ( w8499 , w8498 );
and ( w8500 , w8499 , w8326 );
and ( w8501 , w8500 , w8281 );
and ( w8502 , w8501 , g2 );
nor ( w8503 , w8502 , w7824 );
and ( w8504 , w8503 , g13 );
and ( w8505 , w8504 , g11 );
nor ( w8506 , w8505 , w8448 );
not ( w8507 , w8506 );
and ( w8508 , w8507 , w8491 );
nor ( w8509 , w8373 , w8508 );
not ( w8510 , w8509 );
and ( w8511 , w8510 , w213 );
not ( w8512 , w8511 );
and ( w8513 , w8512 , w8326 );
and ( w8514 , w8513 , w8281 );
and ( w8515 , w8514 , g2 );
nor ( w8516 , w8515 , w7824 );
and ( w8517 , w8516 , g13 );
not ( w8518 , w8517 );
and ( w8519 , w8347 , w8518 );
and ( w8520 , w8519 , w4357 );
not ( w8521 , w8520 );
and ( w8522 , w8521 , w8366 );
not ( w8523 , w8522 );
and ( w8524 , w8523 , g6 );
not ( w8525 , w8524 );
and ( w8526 , w8525 , w8115 );
and ( w8527 , w8526 , w8837 );
and ( w8528 , w8527 , g16 );
nor ( w8529 , w8528 , w8508 );
not ( w8530 , w8529 );
and ( w8531 , w8530 , w213 );
nor ( w8532 , w8531 , g1 );
not ( w8533 , w8532 );
and ( w8534 , w8533 , g14 );
not ( w8535 , w8534 );
and ( w8536 , w8535 , w8326 );
and ( w8537 , w8536 , w8281 );
and ( w8538 , w8537 , g2 );
nor ( w8539 , w8538 , w7824 );
and ( w8540 , w8539 , g13 );
nor ( w8541 , w8068 , w8540 );
not ( w8542 , w8541 );
and ( w8543 , w8542 , g16 );
nor ( w8544 , w8543 , w8508 );
not ( w8545 , w8544 );
and ( w8546 , w8545 , w213 );
nor ( w8547 , w8546 , g1 );
and ( w8548 , w8547 , w8326 );
and ( w8549 , w8548 , w8281 );
and ( w8550 , w8549 , g2 );
nor ( w8551 , w8550 , w7824 );
and ( w8552 , w8551 , g13 );
not ( w8553 , w1516 );
and ( w8554 , w8553 , w8552 );
nor ( w8555 , w8554 , w8540 );
and ( w8556 , w8555 , w8792 );
and ( w8557 , w8556 , w8281 );
and ( w8558 , w8557 , g2 );
nor ( w8559 , w8558 , w7824 );
not ( w8560 , w7835 );
and ( w8561 , w8560 , w8559 );
not ( w8562 , w8561 );
and ( w8563 , w8562 , g2 );
nor ( w8564 , w8563 , w7824 );
and ( w8565 , g1 , w8860 );
and ( w8566 , w8565 , g3 );
nor ( w8567 , w8566 , g4 );
not ( w8568 , w8567 );
and ( w8569 , w8568 , g12 );
nor ( w8570 , w8569 , g11 );
not ( w8571 , w8570 );
and ( w8572 , w8571 , w4849 );
nor ( w8573 , w8572 , g16 );
not ( w8574 , w8573 );
and ( w8575 , w8574 , g1 );
not ( w8576 , w8575 );
and ( w8577 , w8576 , g13 );
not ( w8578 , w8577 );
and ( w8579 , w8578 , w2585 );
not ( w8580 , w8579 );
and ( w8581 , w8580 , w8062 );
not ( w8582 , w8581 );
and ( w8583 , w8582 , g1 );
and ( w8584 , w5802 , w8828 );
and ( w8585 , w8584 , w8837 );
nor ( w8586 , w8585 , g1 );
not ( w8587 , w8586 );
and ( w8588 , w8587 , g13 );
not ( w8589 , w8588 );
and ( w8590 , w8589 , g2 );
and ( w8591 , w8590 , g6 );
not ( w8592 , w8591 );
and ( w8593 , w8592 , g6 );
nor ( w8594 , w8593 , g1 );
and ( w8595 , w8594 , g2 );
nor ( w8596 , w8583 , w8595 );
not ( w8597 , w3601 );
and ( w8598 , w8597 , w8062 );
and ( w8599 , w8598 , w8559 );
and ( w8600 , w8599 , w213 );
not ( w8601 , w8600 );
and ( w8602 , w8601 , w8326 );
not ( w8603 , w8596 );
and ( w8604 , w8603 , w8602 );
and ( w8605 , w8604 , g2 );
nor ( w8606 , w8605 , w7824 );
and ( w8607 , w8606 , g13 );
nor ( w8608 , w8564 , w8607 );
not ( w8609 , w8608 );
and ( w8610 , w8609 , g16 );
nor ( w8611 , w7826 , w8606 );
and ( w8612 , w8611 , w4912 );
nor ( w8613 , w8612 , w8608 );
not ( w8614 , w8613 );
and ( w8615 , w8614 , g2 );
nor ( w8616 , w8615 , g16 );
and ( w8617 , w8616 , w8559 );
and ( w8618 , w8617 , w8819 );
nor ( w8619 , w8618 , w8607 );
not ( w8620 , w8610 );
and ( w8621 , w8620 , w8619 );
nor ( w8622 , w8621 , g13 );
nor ( w8623 , w8622 , w8607 );
and ( w8624 , w7833 , w8623 );
and ( w8625 , w8624 , w8833 );
and ( w8626 , w8625 , g1 );
not ( w8627 , w8626 );
and ( w8628 , w8627 , w8559 );
and ( w8629 , w8628 , w8819 );
nor ( w8630 , w8629 , w8607 );
nor ( w8631 , w7829 , w8630 );
not ( w8632 , w8631 );
and ( w8633 , w8632 , g1 );
and ( w8634 , w8633 , g8 );
not ( w8635 , w8634 );
and ( w8636 , w8635 , g8 );
not ( w8637 , w8636 );
and ( w8638 , w8637 , w7040 );
and ( w8639 , w8638 , w8845 );
and ( w8640 , w8639 , w400 );
and ( w8641 , w8640 , w8828 );
and ( w8642 , w8641 , g11 );
and ( w8643 , w8642 , w8623 );
not ( w8644 , w8643 );
and ( w8645 , w8644 , w8559 );
and ( w8646 , w8645 , w8819 );
nor ( w8647 , w8646 , w8607 );
and ( w8648 , w8647 , w8828 );
and ( w8649 , w8648 , g9 );
and ( w8650 , w8608 , w8765 );
and ( w8651 , w8650 , g16 );
and ( w8652 , w8651 , w8833 );
and ( w8653 , w8652 , g1 );
not ( w8654 , w8653 );
and ( w8655 , w8654 , w8559 );
and ( w8656 , w8655 , w8819 );
nor ( w8657 , w8656 , w8607 );
nor ( w8658 , w8649 , w8657 );
not ( w8659 , w8658 );
and ( w8660 , w8659 , g11 );
not ( w8661 , w8660 );
and ( w8662 , w8661 , g14 );
not ( w8663 , w8662 );
and ( w8664 , w8663 , w8623 );
not ( w8665 , w8664 );
and ( w8666 , w8665 , w8559 );
and ( w8667 , w8666 , w8819 );
nor ( w8668 , w8667 , w8607 );
nor ( w8669 , w8668 , w8657 );
nor ( w8670 , w8669 , g9 );
nor ( w8671 , w8670 , g13 );
and ( w8672 , w4449 , w8831 );
not ( w8673 , w8672 );
and ( w8674 , w8673 , g9 );
nor ( w8675 , w8674 , w8669 );
nor ( w8676 , w1430 , w8669 );
and ( w8677 , w8675 , w8676 );
and ( w8678 , w8677 , g3 );
and ( w8679 , w8678 , g17 );
and ( w8680 , w8679 , w4849 );
not ( w8681 , w8680 );
and ( w8682 , w8681 , g13 );
not ( w8683 , w8682 );
and ( w8684 , w8683 , g1 );
and ( w8685 , w8684 , g6 );
not ( w8686 , w8685 );
and ( w8687 , w8686 , g11 );
nor ( w8688 , w8671 , w8687 );
and ( w8689 , w8688 , g1 );
and ( w8690 , w1517 , w8831 );
nor ( w8691 , w8669 , w7826 );
and ( w8692 , w8691 , g9 );
and ( w8693 , w8692 , w4912 );
nor ( w8694 , w8693 , w8670 );
nor ( w8695 , w8694 , g6 );
and ( w8696 , w8695 , w7040 );
and ( w8697 , w8696 , g1 );
nor ( w8698 , w7905 , w8607 );
and ( w8699 , w8698 , w8845 );
and ( w8700 , w8699 , g2 );
nor ( w8701 , g1 , w8698 );
nor ( w8702 , w8701 , g6 );
and ( w8703 , w8702 , w8831 );
nor ( w8704 , w8690 , w8703 );
not ( w8705 , w8704 );
and ( w8706 , w8705 , g3 );
and ( w8707 , w1517 , w8730 );
and ( w8708 , w8707 , w8735 );
nor ( w8709 , w8708 , w33 );
not ( w8710 , w3188 );
and ( w8711 , w8710 , g6 );
not ( w8712 , w8709 );
and ( w8713 , w8712 , w8711 );
and ( w8714 , w8713 , w8831 );
nor ( w8715 , g3 , w8669 );
and ( w8716 , w8714 , w8715 );
and ( w8717 , w8716 , g2 );
and ( w8718 , w8715 , w8845 );
nor ( w8719 , w8717 , w8718 );
not ( w8720 , w8717 );
and ( w8721 , g6 , w8720 );
and ( w8722 , w8721 , w8735 );
nor ( w8723 , w8722 , g1 );
not ( w8724 , w8719 );
and ( w8725 , w8724 , w8723 );
and ( w8726 , w8725 , g4 );
nor ( w8727 , g14 , g9 );
not ( w8728 , g12 );
and ( w8729 , w8727 , w8728 );
not ( w8730 , g10 );
and ( w8731 , w8729 , w8730 );
and ( w8732 , w8731 , w8819 );
and ( w8733 , w8732 , w8845 );
and ( w8734 , w8733 , g15 );
not ( w8735 , g3 );
and ( w8736 , w8735 , w8734 );
nor ( w8737 , w8700 , g6 );
nor ( w8738 , w8737 , w8669 );
and ( w8739 , w19 , w33 );
nor ( w8740 , w8739 , g5 );
and ( w8741 , w8740 , g10 );
not ( w8742 , g7 );
and ( w8743 , w8741 , w8742 );
nor ( w8744 , w8743 , g8 );
nor ( w8745 , w8744 , g8 );
nor ( w8746 , w8745 , g9 );
and ( w8747 , w8746 , w8831 );
and ( w8748 , w6484 , g10 );
not ( w8749 , w8748 );
and ( w8750 , w8749 , w1244 );
nor ( w8751 , w8750 , g7 );
nor ( w8752 , w8751 , g1 );
and ( w8753 , w8752 , w8767 );
nor ( w8754 , w8753 , g8 );
not ( w8755 , w8754 );
and ( w8756 , w8755 , g6 );
and ( w8757 , w8756 , w8831 );
and ( w8758 , w8747 , w8757 );
and ( w8759 , w8758 , w361 );
and ( w8760 , w8759 , w408 );
and ( w8761 , w8760 , w27 );
nor ( w8762 , w8672 , w8761 );
and ( w8763 , w2177 , w8767 );
nor ( w8764 , w8763 , g7 );
not ( w8765 , g9 );
and ( w8766 , w8764 , w8765 );
not ( w8767 , g8 );
and ( w8768 , w8766 , w8767 );
not ( w8769 , g5 );
and ( w8770 , w8768 , w8769 );
nor ( w8771 , w8770 , g1 );
and ( w8772 , w8771 , w8831 );
not ( w8773 , w8762 );
and ( w8774 , w8773 , w8772 );
and ( w8775 , w8774 , g2 );
and ( w8776 , w5579 , w8831 );
and ( w8777 , w8776 , w8845 );
nor ( w8778 , w8775 , w8777 );
nor ( w8779 , w8778 , g3 );
not ( w8780 , w8734 );
and ( w8781 , w8779 , w8780 );
and ( w8782 , w8781 , w27 );
not ( w8783 , w8782 );
and ( w8784 , w8783 , g16 );
not ( w8785 , w8784 );
and ( w8786 , w8785 , w8776 );
nor ( w8787 , w8786 , g11 );
not ( w8788 , w8787 );
and ( w8789 , w8788 , g2 );
and ( w8790 , w8738 , w8789 );
and ( w8791 , w8738 , g3 );
not ( w8792 , g1 );
and ( w8793 , w8791 , w8792 );
and ( w8794 , w8793 , g2 );
nor ( w8795 , w8790 , w8794 );
not ( w8796 , w8795 );
and ( w8797 , w8796 , w8776 );
not ( w8798 , w8736 );
and ( w8799 , w8798 , w8797 );
not ( w8800 , w8799 );
and ( w8801 , w8800 , g16 );
not ( w8802 , w8801 );
and ( w8803 , w8802 , w8776 );
nor ( w8804 , w8803 , g11 );
not ( w8805 , w8804 );
and ( w8806 , w8805 , g2 );
nor ( w8807 , w8726 , w8806 );
nor ( w8808 , w8807 , g1 );
and ( w8809 , w8808 , g2 );
nor ( w8810 , w8706 , w8809 );
not ( w8811 , w8810 );
and ( w8812 , w8811 , w8723 );
and ( w8813 , w8812 , g4 );
nor ( w8814 , w8813 , w8806 );
nor ( w8815 , w8814 , g1 );
and ( w8816 , w8815 , g2 );
and ( w8817 , w8700 , w8816 );
nor ( w8818 , w8697 , w8817 );
not ( w8819 , g13 );
and ( w8820 , w8818 , w8819 );
not ( w8821 , w8817 );
and ( w8822 , w8821 , g13 );
and ( w8823 , w8822 , w8828 );
and ( w8824 , w8823 , g11 );
and ( w8825 , w4803 , g6 );
and ( w8826 , w8825 , g13 );
and ( w8827 , w8826 , g10 );
not ( w8828 , g16 );
and ( w8829 , w8827 , w8828 );
nor ( w8830 , w3004 , w8829 );
not ( w8831 , w8669 );
and ( w8832 , w8830 , w8831 );
not ( w8833 , g15 );
and ( w8834 , w8832 , w8833 );
and ( w8835 , w8834 , g1 );
nor ( w8836 , w8835 , w8816 );
not ( w8837 , g11 );
and ( w8838 , w8836 , w8837 );
not ( w8839 , w8838 );
and ( w8840 , w8839 , g2 );
not ( w8841 , w8824 );
and ( w8842 , w8841 , w8840 );
not ( w8843 , w8820 );
and ( w8844 , w8843 , w8842 );
not ( w8845 , g6 );
and ( w8846 , w8844 , w8845 );
and ( w8847 , w1517 , w8840 );
not ( w8848 , w8847 );
and ( w8849 , w1588 , w8848 );
not ( w8850 , w8849 );
and ( w8851 , w8850 , g2 );
and ( w8852 , w8851 , g6 );
and ( w8853 , w27 , g2 );
nor ( w8854 , w8853 , g3 );
nor ( w8855 , w8854 , g9 );
nor ( w8856 , w8855 , g9 );
nor ( w8857 , w8856 , g1 );
not ( w8858 , w8857 );
and ( w8859 , w8858 , g15 );
not ( w8860 , g4 );
and ( w8861 , w8859 , w8860 );
nor ( w8862 , w8861 , g6 );
and ( w8863 , w8862 , w8840 );
nor ( w8864 , w8852 , w8863 );
nor ( w8865 , w8864 , w8669 );
and ( w8866 , w8865 , w8840 );
and ( w8867 , w8846 , w8866 );
nor ( w8868 , w8867 , g16 );
and ( w8869 , w8868 , g11 );
not ( w8870 , w8869 );
and ( w8871 , w8870 , w8840 );
nor ( w8872 , w8690 , w8871 );
not ( w8873 , w8872 );
and ( w8874 , w8873 , w8866 );
nor ( w8875 , w8689 , w8874 );
not ( w8876 , w8875 );
and ( w8877 , w8876 , g2 );
and ( w8878 , w8877 , g6 );
nor ( w8879 , w8878 , w8871 );
not ( w8880 , w8879 );
and ( w8881 , w8880 , w8866 );
nor ( t_11 , w7824 , w8881 );

endmodule
