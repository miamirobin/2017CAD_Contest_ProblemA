module patch (t_0, g1, g2, g3);
input g1, g2, g3;
output t_0;
wire w1, w2, w3, w4, w5, w6;

not ( w1 , g1 );
and ( w2 , w1 , g2 );
and ( w3 , g1 , g3 );
nor ( w4 , g1 , g3 );
nor ( w5 , w3 , w4 );
nor ( w6 , w5 , g2 );
nor ( t_0 , w2 , w6 );

endmodule
