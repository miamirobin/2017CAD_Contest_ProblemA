module patch (t_0, t_1, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13;
output t_0, t_1;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572;

and ( w1 , g1 , w202 );
not ( w2 , w1 );
and ( w3 , w2 , g3 );
and ( w4 , g1 , g4 );
and ( w5 , w3 , w4 );
and ( w6 , w5 , g1 );
and ( w7 , w224 , g4 );
nor ( w8 , w6 , w7 );
and ( w9 , w202 , g3 );
nor ( w10 , w9 , g2 );
nor ( w11 , w8 , w10 );
and ( w12 , w11 , g3 );
and ( w13 , g5 , g1 );
and ( w14 , w3 , w13 );
not ( w15 , w14 );
and ( w16 , w15 , g1 );
not ( w17 , w16 );
and ( w18 , w12 , w17 );
and ( w19 , w18 , g1 );
and ( w20 , w224 , g2 );
and ( w21 , w19 , w151 );
and ( w22 , w535 , g7 );
and ( w23 , w22 , w552 );
not ( w24 , w23 );
and ( w25 , w24 , g7 );
and ( w26 , w25 , w552 );
and ( w27 , w26 , w535 );
and ( w28 , g6 , w543 );
and ( w29 , w28 , g9 );
nor ( w30 , w29 , g9 );
nor ( w31 , g9 , w30 );
nor ( w32 , w27 , w31 );
not ( w33 , w21 );
and ( w34 , w33 , w32 );
not ( w35 , w34 );
and ( w36 , w35 , g2 );
and ( w37 , w36 , g10 );
and ( w38 , g8 , w535 );
nor ( w39 , w38 , g6 );
nor ( w40 , w39 , g11 );
not ( w41 , w40 );
and ( w42 , w41 , g8 );
and ( w43 , g7 , w491 );
not ( w44 , w42 );
and ( w45 , w44 , w43 );
not ( w46 , w45 );
and ( w47 , w46 , g7 );
nor ( w48 , w47 , g9 );
and ( w49 , w48 , w497 );
and ( w50 , g7 , g6 );
nor ( w51 , w50 , w38 );
not ( w52 , w51 );
and ( w53 , w52 , g8 );
not ( w54 , w53 );
and ( w55 , w54 , g8 );
nor ( w56 , g12 , g9 );
not ( w57 , w55 );
and ( w58 , w57 , w56 );
nor ( w59 , w58 , g12 );
not ( w60 , w59 );
and ( w61 , w60 , g7 );
and ( w62 , w49 , w61 );
and ( w63 , w62 , w497 );
nor ( w64 , w63 , g11 );
not ( w65 , w64 );
and ( w66 , w65 , w43 );
and ( w67 , w66 , g7 );
nor ( w68 , g9 , w67 );
not ( w69 , w68 );
and ( w70 , w69 , g7 );
and ( w71 , w70 , g13 );
not ( w72 , w71 );
and ( w73 , w72 , w70 );
not ( w74 , w73 );
and ( w75 , w74 , g13 );
not ( w76 , w75 );
and ( w77 , w76 , g13 );
nor ( w78 , w77 , g5 );
and ( w79 , w78 , w202 );
and ( w80 , w79 , w224 );
and ( w81 , w80 , g4 );
not ( w82 , w81 );
and ( w83 , w82 , w32 );
not ( w84 , w83 );
and ( w85 , w84 , g3 );
not ( w86 , w77 );
and ( w87 , w86 , g1 );
and ( w88 , w87 , w219 );
and ( w89 , w88 , g2 );
and ( w90 , w89 , g5 );
not ( w91 , w90 );
and ( w92 , w91 , w32 );
nor ( w93 , w92 , g3 );
not ( w94 , w93 );
and ( w95 , w94 , w32 );
not ( w96 , w95 );
and ( w97 , w96 , g10 );
not ( w98 , w97 );
and ( w99 , w98 , w32 );
not ( w100 , w85 );
and ( w101 , w100 , w99 );
not ( w102 , w101 );
and ( w103 , w102 , g10 );
nor ( w104 , w77 , g3 );
and ( w105 , w104 , g1 );
and ( w106 , w105 , w232 );
not ( w107 , w106 );
and ( w108 , w107 , g1 );
nor ( w109 , w108 , g10 );
and ( w110 , w109 , g2 );
and ( w111 , w4 , g2 );
and ( w112 , w111 , w228 );
and ( w113 , w110 , w112 );
nor ( w114 , g2 , g1 );
nor ( w115 , w114 , w13 );
not ( w116 , w115 );
and ( w117 , w116 , g4 );
not ( w118 , w13 );
and ( w119 , g1 , w118 );
not ( w120 , w119 );
and ( w121 , w120 , w3 );
and ( w122 , w117 , w121 );
nor ( w123 , w113 , w122 );
nor ( w124 , w123 , g10 );
nor ( w125 , w103 , w124 );
and ( w126 , w149 , g3 );
and ( w127 , w126 , g2 );
and ( w128 , w127 , g5 );
not ( w129 , w128 );
and ( w130 , w129 , g2 );
and ( w131 , w130 , g5 );
not ( w132 , w131 );
and ( w133 , w132 , w3 );
and ( w134 , w133 , w4 );
nor ( w135 , w134 , w7 );
and ( w136 , g5 , g3 );
and ( w137 , w136 , w202 );
nor ( w138 , w137 , g2 );
nor ( w139 , w135 , w138 );
not ( w140 , w114 );
and ( w141 , w139 , w140 );
not ( w142 , w138 );
and ( w143 , w142 , w7 );
and ( w144 , w143 , w18 );
and ( w145 , w144 , w149 );
nor ( w146 , w141 , w145 );
nor ( w147 , w146 , w16 );
and ( w148 , w147 , g3 );
not ( w149 , g10 );
and ( w150 , w148 , w149 );
not ( w151 , w20 );
and ( w152 , w150 , w151 );
nor ( w153 , w152 , w112 );
nor ( w154 , w150 , w112 );
nor ( w155 , w154 , g10 );
not ( w156 , w153 );
and ( w157 , w156 , w155 );
and ( w158 , w552 , w28 );
not ( w159 , w158 );
and ( w160 , w159 , g6 );
and ( w161 , w160 , w543 );
and ( w162 , g12 , g9 );
not ( w163 , w161 );
and ( w164 , w163 , w162 );
nor ( w165 , w164 , g8 );
and ( w166 , w165 , g12 );
and ( w167 , w166 , g9 );
nor ( w168 , w77 , w167 );
and ( w169 , w168 , g10 );
and ( w170 , w169 , w232 );
and ( w171 , w170 , g3 );
and ( w172 , w171 , w202 );
and ( w173 , w172 , w7 );
and ( w174 , g1 , w219 );
and ( w175 , w174 , g2 );
not ( w176 , w175 );
and ( w177 , w176 , w32 );
nor ( w178 , w177 , g3 );
and ( w179 , w178 , g5 );
nor ( w180 , g2 , g4 );
and ( w181 , w180 , w232 );
nor ( w182 , w179 , w181 );
not ( w183 , w182 );
and ( w184 , w183 , g10 );
and ( w185 , w184 , w228 );
nor ( w186 , w173 , w185 );
not ( w187 , w157 );
and ( w188 , w187 , w186 );
nor ( w189 , w125 , w188 );
nor ( w190 , w37 , w189 );
not ( w191 , w190 );
and ( w192 , w191 , g10 );
nor ( w193 , w169 , g5 );
and ( w194 , g2 , g4 );
and ( w195 , w193 , w194 );
and ( w196 , w195 , w7 );
nor ( w197 , w122 , w196 );
not ( w198 , w126 );
and ( w199 , w198 , g3 );
nor ( w200 , w197 , w199 );
and ( w201 , w200 , w126 );
not ( w202 , g2 );
and ( w203 , w168 , w202 );
nor ( w204 , w203 , g2 );
not ( w205 , w204 );
and ( w206 , w205 , w181 );
and ( w207 , w206 , w232 );
nor ( w208 , w207 , g5 );
nor ( w209 , g1 , g4 );
not ( w210 , w208 );
and ( w211 , w210 , w209 );
and ( w212 , w169 , g1 );
and ( w213 , w212 , g2 );
nor ( w214 , w213 , w209 );
not ( w215 , w214 );
and ( w216 , w215 , g5 );
and ( w217 , w228 , g10 );
and ( w218 , w216 , w217 );
not ( w219 , g4 );
and ( w220 , w218 , w219 );
nor ( w221 , w211 , w220 );
not ( w222 , w221 );
and ( w223 , w222 , g10 );
not ( w224 , g1 );
and ( w225 , w224 , g5 );
not ( w226 , w225 );
and ( w227 , w223 , w226 );
not ( w228 , g3 );
and ( w229 , w227 , w228 );
and ( w230 , w229 , w209 );
and ( w231 , w127 , w7 );
not ( w232 , g5 );
and ( w233 , w231 , w232 );
nor ( w234 , w233 , w122 );
not ( w235 , w113 );
and ( w236 , w234 , w235 );
nor ( w237 , w236 , g10 );
nor ( w238 , w230 , w237 );
nor ( w239 , w188 , w238 );
nor ( w240 , w189 , w239 );
not ( w241 , w201 );
and ( w242 , w241 , w240 );
not ( w243 , w192 );
and ( t_0 , w243 , w242 );
and ( w244 , g8 , g6 );
and ( w245 , w244 , w75 );
and ( w246 , w245 , g9 );
and ( w247 , g12 , w75 );
not ( w248 , w247 );
and ( w249 , w248 , g12 );
and ( w250 , g8 , w50 );
nor ( w251 , w250 , w22 );
not ( w252 , w251 );
and ( w253 , w252 , g8 );
and ( w254 , w253 , w491 );
and ( w255 , w254 , g7 );
and ( w256 , w255 , g8 );
and ( w257 , w256 , w491 );
and ( w258 , w257 , w56 );
not ( w259 , w249 );
and ( w260 , w259 , w258 );
and ( w261 , w260 , w491 );
and ( w262 , w261 , g8 );
nor ( w263 , w246 , w262 );
not ( w264 , w263 );
and ( w265 , w264 , g6 );
not ( w266 , w50 );
and ( w267 , w266 , g6 );
nor ( w268 , w267 , g8 );
nor ( w269 , w268 , g8 );
and ( w270 , w405 , g11 );
and ( w271 , g12 , w497 );
nor ( w272 , w270 , w271 );
not ( w273 , w272 );
and ( w274 , w273 , g12 );
and ( w275 , w274 , w491 );
not ( w276 , w275 );
and ( w277 , w276 , g12 );
and ( w278 , w70 , g11 );
not ( w279 , w278 );
and ( w280 , w279 , g11 );
nor ( w281 , g8 , g9 );
and ( w282 , w280 , w281 );
and ( w283 , w23 , g12 );
nor ( w284 , w283 , w280 );
not ( w285 , w284 );
and ( w286 , w285 , w281 );
nor ( w287 , w286 , g9 );
nor ( w288 , g8 , g6 );
not ( w289 , w287 );
and ( w290 , w289 , w288 );
nor ( w291 , w282 , w290 );
nor ( w292 , w283 , g8 );
and ( w293 , w292 , w535 );
and ( w294 , w293 , g9 );
nor ( w295 , w291 , w294 );
not ( w296 , w277 );
and ( w297 , w296 , w295 );
and ( w298 , w297 , g7 );
and ( w299 , w298 , w491 );
and ( w300 , w299 , g13 );
nor ( w301 , g8 , w300 );
not ( w302 , w301 );
and ( w303 , w302 , g7 );
nor ( w304 , w303 , w280 );
nor ( w305 , w304 , g9 );
and ( w306 , w305 , g13 );
nor ( w307 , w306 , g9 );
and ( w308 , w43 , w497 );
and ( w309 , w308 , w38 );
not ( w310 , w307 );
and ( w311 , w310 , w309 );
nor ( w312 , g8 , w295 );
not ( w313 , w312 );
and ( w314 , w313 , g13 );
and ( w315 , w314 , g9 );
and ( w316 , w315 , w485 );
and ( w317 , w316 , g11 );
and ( w318 , w317 , g6 );
nor ( w319 , w318 , w309 );
nor ( w320 , w319 , g7 );
and ( w321 , w320 , g8 );
nor ( w322 , w311 , w321 );
and ( w323 , g7 , w295 );
and ( w324 , w491 , w280 );
nor ( w325 , w324 , g9 );
not ( w326 , w325 );
and ( w327 , w326 , g11 );
not ( w328 , w327 );
and ( w329 , w328 , g11 );
not ( w330 , w329 );
and ( w331 , w330 , w295 );
and ( w332 , w331 , w543 );
and ( w333 , w332 , w552 );
and ( w334 , w333 , g13 );
nor ( w335 , w323 , w334 );
nor ( w336 , w335 , g11 );
nor ( w337 , w336 , g11 );
not ( w338 , w337 );
and ( w339 , w338 , g13 );
not ( w340 , w339 );
and ( w341 , w322 , w340 );
not ( w342 , w265 );
and ( w343 , w342 , w341 );
and ( w344 , g12 , w244 );
nor ( w345 , w344 , w309 );
not ( w346 , w345 );
and ( w347 , w346 , g9 );
and ( w348 , w497 , w314 );
and ( w349 , w348 , g6 );
and ( w350 , w309 , w535 );
and ( w351 , w350 , g8 );
nor ( w352 , w349 , w351 );
nor ( w353 , w352 , g9 );
and ( w354 , w353 , g7 );
nor ( w355 , w354 , w321 );
not ( w356 , w347 );
and ( w357 , w356 , w355 );
not ( w358 , w357 );
and ( w359 , w358 , g7 );
nor ( w360 , w359 , w321 );
not ( w361 , w335 );
and ( w362 , w361 , g13 );
not ( w363 , w362 );
and ( w364 , w360 , w363 );
not ( w365 , w364 );
and ( w366 , w365 , g13 );
not ( w367 , w343 );
and ( w368 , w367 , w366 );
and ( w369 , g13 , g11 );
and ( w370 , w368 , w369 );
nor ( w371 , w267 , g9 );
and ( w372 , w371 , g12 );
not ( w373 , g13 );
and ( w374 , w372 , w373 );
and ( w375 , w374 , w497 );
nor ( w376 , w375 , g13 );
and ( w377 , w247 , w268 );
and ( w378 , w377 , g6 );
nor ( w379 , w378 , w22 );
nor ( w380 , w379 , g8 );
and ( w381 , w380 , w491 );
and ( w382 , w381 , g13 );
not ( w383 , w382 );
and ( w384 , w383 , g13 );
nor ( w385 , w384 , g11 );
and ( w386 , w385 , w271 );
and ( w387 , w386 , w491 );
and ( w388 , g7 , w552 );
and ( w389 , w387 , w388 );
and ( w390 , w389 , w552 );
not ( w391 , w376 );
and ( w392 , w391 , w390 );
and ( w393 , w392 , w497 );
not ( w394 , w369 );
and ( w395 , w394 , g13 );
not ( w396 , w70 );
and ( w397 , w396 , g7 );
nor ( w398 , w395 , w397 );
and ( w399 , w398 , w491 );
and ( w400 , w552 , g6 );
and ( w401 , w399 , w400 );
not ( w402 , w401 );
and ( w403 , w402 , g6 );
nor ( w404 , w403 , g9 );
not ( w405 , w269 );
and ( w406 , w404 , w405 );
and ( w407 , g12 , g11 );
and ( w408 , w406 , w407 );
and ( w409 , w408 , g7 );
not ( w410 , w409 );
and ( w411 , w410 , g7 );
nor ( w412 , w411 , g8 );
nor ( w413 , w412 , g8 );
nor ( w414 , w413 , g9 );
nor ( w415 , w393 , w414 );
not ( w416 , w415 );
and ( w417 , w416 , g12 );
and ( w418 , w267 , g7 );
not ( w419 , w418 );
and ( w420 , w419 , g8 );
not ( w421 , w420 );
and ( w422 , w421 , g13 );
not ( w423 , w422 );
and ( w424 , w423 , g13 );
nor ( w425 , w424 , g12 );
nor ( w426 , g12 , g11 );
and ( w427 , w425 , w426 );
nor ( w428 , w427 , g11 );
nor ( w429 , w428 , g12 );
and ( w430 , w429 , w56 );
and ( w431 , w430 , w43 );
and ( w432 , w431 , w388 );
not ( w433 , w432 );
and ( w434 , w433 , g7 );
nor ( w435 , w434 , g8 );
and ( w436 , w435 , w491 );
nor ( w437 , w436 , g9 );
not ( w438 , w417 );
and ( w439 , w438 , w437 );
and ( w440 , w439 , w497 );
and ( w441 , w440 , g7 );
and ( w442 , w441 , g6 );
nor ( w443 , w442 , g12 );
and ( w444 , w443 , w491 );
not ( w445 , w444 );
and ( w446 , w445 , g7 );
and ( w447 , w446 , g8 );
and ( w448 , w295 , w497 );
and ( w449 , w448 , w552 );
nor ( w450 , w447 , w449 );
nor ( w451 , w450 , g11 );
and ( w452 , w451 , g13 );
nor ( w453 , w370 , w452 );
nor ( w454 , w442 , w311 );
not ( w455 , w454 );
and ( w456 , w455 , g13 );
and ( w457 , w485 , g9 );
and ( w458 , w280 , w457 );
and ( w459 , w458 , g13 );
nor ( w460 , g7 , w459 );
not ( w461 , w460 );
and ( w462 , w461 , w244 );
nor ( w463 , w462 , w309 );
not ( w464 , w463 );
and ( w465 , w464 , g9 );
and ( w466 , w465 , g13 );
nor ( w467 , w456 , w466 );
not ( w468 , w467 );
and ( w469 , w468 , g11 );
nor ( w470 , w288 , w244 );
not ( w471 , w470 );
and ( w472 , w471 , g7 );
and ( w473 , w472 , g12 );
and ( w474 , w244 , w543 );
and ( w475 , w474 , g11 );
and ( w476 , w475 , w485 );
and ( w477 , w476 , g13 );
nor ( w478 , w473 , w477 );
not ( w479 , w478 );
and ( w480 , w479 , g9 );
and ( w481 , w22 , w497 );
and ( w482 , w481 , g12 );
and ( w483 , w497 , g6 );
and ( w484 , w483 , g7 );
not ( w485 , g12 );
and ( w486 , w484 , w485 );
and ( w487 , w486 , w491 );
nor ( w488 , w482 , w487 );
not ( w489 , w488 );
and ( w490 , w489 , g8 );
not ( w491 , g9 );
and ( w492 , w490 , w491 );
and ( w493 , w492 , g13 );
nor ( w494 , w480 , w493 );
not ( w495 , w494 );
and ( w496 , w495 , g13 );
not ( w497 , g11 );
and ( w498 , w496 , w497 );
nor ( w499 , w469 , w498 );
not ( w500 , w499 );
and ( w501 , w500 , g6 );
nor ( w502 , w501 , w309 );
nor ( w503 , g11 , g6 );
and ( w504 , w503 , w552 );
not ( w505 , w504 );
and ( w506 , w502 , w505 );
not ( w507 , w506 );
and ( w508 , w507 , g12 );
and ( w509 , w508 , g9 );
not ( w510 , w407 );
and ( w511 , w510 , g12 );
not ( w512 , w511 );
and ( w513 , w512 , g9 );
not ( w514 , w513 );
and ( w515 , w514 , g11 );
and ( w516 , w515 , w535 );
nor ( w517 , w516 , g6 );
not ( w518 , w517 );
and ( w519 , w518 , g12 );
not ( w520 , w519 );
and ( w521 , w520 , g12 );
not ( w522 , w521 );
and ( w523 , w522 , w295 );
and ( w524 , w523 , g13 );
nor ( w525 , w456 , w524 );
not ( w526 , w509 );
and ( w527 , w526 , w525 );
and ( w528 , g6 , w295 );
not ( w529 , w528 );
and ( w530 , w529 , g6 );
not ( w531 , w530 );
and ( w532 , w531 , g7 );
not ( w533 , w532 );
and ( w534 , w533 , g7 );
not ( w535 , g6 );
and ( w536 , w535 , g12 );
and ( w537 , w536 , g9 );
and ( w538 , w537 , g7 );
and ( w539 , w538 , g11 );
nor ( w540 , w539 , g8 );
nor ( w541 , w540 , g8 );
nor ( w542 , w534 , w541 );
not ( w543 , g7 );
and ( w544 , w295 , w543 );
nor ( w545 , w544 , g7 );
not ( w546 , w545 );
and ( w547 , w546 , g9 );
not ( w548 , w547 );
and ( w549 , w548 , g9 );
not ( w550 , w549 );
and ( w551 , w542 , w550 );
not ( w552 , g8 );
and ( w553 , w551 , w552 );
nor ( w554 , w553 , g8 );
not ( w555 , w554 );
and ( w556 , w555 , g13 );
not ( w557 , w527 );
and ( w558 , w557 , w556 );
and ( w559 , w558 , g7 );
not ( w560 , w162 );
and ( w561 , w560 , g12 );
not ( w562 , w561 );
and ( w563 , w562 , g11 );
not ( w564 , w563 );
and ( w565 , w564 , g11 );
not ( w566 , w565 );
and ( w567 , w566 , w295 );
and ( w568 , w567 , g13 );
not ( w569 , w568 );
and ( w570 , w319 , w569 );
nor ( w571 , w570 , g7 );
nor ( w572 , w559 , w571 );
or ( t_1 , w453 , w572 );

endmodule
