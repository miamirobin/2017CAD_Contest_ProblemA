module patch (t_0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13;
output t_0;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202;

and ( w1 , g2 , w110 );
nor ( w2 , g1 , w1 );
not ( w3 , g5 );
and ( w4 , g4 , w3 );
nor ( w5 , w4 , g6 );
not ( w6 , w5 );
and ( w7 , w6 , g7 );
and ( w8 , w7 , w110 );
and ( w9 , w2 , w86 );
not ( w10 , g4 );
and ( w11 , w10 , g5 );
nor ( w12 , w11 , w8 );
and ( w13 , w12 , g7 );
and ( w14 , w13 , w110 );
and ( w15 , w9 , w14 );
nor ( w16 , g4 , g6 );
not ( w17 , w16 );
and ( w18 , w17 , g5 );
nor ( w19 , g4 , g5 );
nor ( w20 , w19 , g3 );
not ( w21 , w20 );
and ( w22 , w21 , g7 );
nor ( w23 , w18 , w22 );
and ( w24 , w23 , w1 );
and ( w25 , g8 , w110 );
nor ( w26 , w24 , w25 );
and ( w27 , w2 , w20 );
not ( w28 , g9 );
and ( w29 , w28 , g10 );
nor ( w30 , w29 , g3 );
not ( w31 , g11 );
and ( w32 , w31 , g3 );
nor ( w33 , w30 , w32 );
and ( w34 , w33 , w106 );
not ( w35 , g10 );
and ( w36 , g9 , w35 );
nor ( w37 , w36 , g12 );
nor ( w38 , w37 , g3 );
nor ( w39 , w38 , g12 );
nor ( w40 , w39 , g11 );
nor ( w41 , w34 , w40 );
and ( w42 , w27 , w41 );
nor ( w43 , w14 , w42 );
and ( w44 , w23 , g7 );
nor ( w45 , w2 , w25 );
and ( w46 , w45 , w151 );
nor ( w47 , g13 , w25 );
nor ( w48 , w47 , w1 );
and ( w49 , w48 , w153 );
nor ( w50 , w46 , w49 );
nor ( w51 , w44 , w50 );
nor ( w52 , w51 , g1 );
and ( w53 , w52 , w181 );
and ( w54 , w25 , w1 );
nor ( w55 , w54 , g13 );
and ( w56 , w55 , w153 );
and ( w57 , g13 , g1 );
nor ( w58 , w57 , w25 );
and ( w59 , w58 , w181 );
nor ( w60 , w56 , w59 );
and ( w61 , w14 , w60 );
nor ( w62 , w53 , w61 );
nor ( w63 , w43 , w62 );
not ( w64 , w63 );
and ( w65 , w64 , w25 );
nor ( w66 , g13 , g1 );
not ( w67 , w66 );
and ( w68 , w67 , w59 );
nor ( w69 , g7 , g6 );
nor ( w70 , w68 , w69 );
and ( w71 , g7 , g6 );
and ( w72 , w70 , w89 );
not ( w73 , g7 );
and ( w74 , w73 , g6 );
and ( w75 , w118 , g1 );
nor ( w76 , w75 , g13 );
nor ( w77 , w20 , g6 );
and ( w78 , w77 , g7 );
nor ( w79 , w78 , w74 );
and ( w80 , w79 , w153 );
not ( w81 , w80 );
and ( w82 , w81 , g13 );
not ( w83 , w82 );
and ( w84 , w83 , w79 );
and ( w85 , w84 , w41 );
not ( w86 , w8 );
and ( w87 , w1 , w86 );
nor ( w88 , w87 , g1 );
not ( w89 , w71 );
and ( w90 , w89 , g1 );
nor ( w91 , w90 , w1 );
and ( w92 , w91 , g3 );
nor ( w93 , w88 , w92 );
nor ( w94 , w93 , w25 );
and ( w95 , w94 , w151 );
and ( w96 , w199 , w25 );
nor ( w97 , g1 , w69 );
not ( w98 , w97 );
and ( w99 , w98 , g13 );
nor ( w100 , g11 , g12 );
and ( w101 , g11 , g12 );
nor ( w102 , w100 , w101 );
nor ( w103 , g10 , g9 );
and ( w104 , g10 , g9 );
nor ( w105 , w104 , g11 );
not ( w106 , g12 );
and ( w107 , w105 , w106 );
not ( w108 , w103 );
and ( w109 , w108 , w107 );
not ( w110 , g3 );
and ( w111 , w109 , w110 );
nor ( w112 , w102 , w111 );
nor ( w113 , w99 , w112 );
not ( w114 , w96 );
and ( w115 , w114 , w113 );
not ( w116 , w95 );
and ( w117 , w116 , w115 );
not ( w118 , w74 );
and ( w119 , w118 , g3 );
nor ( w120 , w68 , w25 );
and ( w121 , w120 , w181 );
and ( w122 , w119 , w121 );
and ( w123 , w2 , w44 );
nor ( w124 , w123 , w25 );
not ( w125 , w124 );
and ( w126 , w23 , w125 );
nor ( w127 , w126 , w41 );
not ( w128 , w127 );
and ( w129 , w128 , g7 );
nor ( w130 , w122 , w129 );
and ( w131 , w130 , w201 );
and ( w132 , w153 , g13 );
not ( w133 , w132 );
and ( w134 , w79 , w133 );
nor ( w135 , w134 , w41 );
not ( w136 , w135 );
and ( w137 , g3 , w136 );
nor ( w138 , w137 , w44 );
nor ( w139 , w131 , w138 );
nor ( w140 , w69 , w71 );
and ( w141 , g1 , w140 );
and ( w142 , w79 , w121 );
nor ( w143 , w141 , w142 );
not ( w144 , w143 );
and ( w145 , w144 , g3 );
nor ( w146 , w145 , w25 );
and ( w147 , w1 , w14 );
not ( w148 , w147 );
and ( w149 , w148 , w124 );
and ( w150 , w146 , w149 );
not ( w151 , g13 );
and ( w152 , w150 , w151 );
not ( w153 , g1 );
and ( w154 , w153 , w140 );
nor ( w155 , w154 , w142 );
not ( w156 , w155 );
and ( w157 , w156 , g3 );
not ( w158 , w157 );
and ( w159 , w158 , g13 );
nor ( w160 , w159 , w25 );
and ( w161 , w160 , w181 );
nor ( w162 , w1 , w14 );
nor ( w163 , w61 , g13 );
not ( w164 , w162 );
and ( w165 , w164 , w163 );
not ( w166 , w165 );
and ( w167 , w166 , w25 );
nor ( w168 , w167 , g13 );
nor ( w169 , w161 , w168 );
nor ( w170 , w152 , w169 );
and ( w171 , w139 , w170 );
not ( w172 , w112 );
and ( w173 , w171 , w172 );
nor ( w174 , w117 , w173 );
not ( w175 , w174 );
and ( w176 , w175 , w170 );
nor ( w177 , w85 , w176 );
nor ( w178 , w76 , w177 );
and ( w179 , w178 , w79 );
nor ( w180 , w179 , w25 );
not ( w181 , w1 );
and ( w182 , w180 , w181 );
not ( w183 , w182 );
and ( w184 , w183 , w41 );
nor ( w185 , w184 , w176 );
not ( w186 , w72 );
and ( w187 , w186 , w185 );
not ( w188 , w187 );
and ( w189 , w188 , w41 );
nor ( w190 , w189 , w176 );
nor ( w191 , w65 , w190 );
and ( w192 , w191 , w41 );
nor ( w193 , w192 , w176 );
nor ( w194 , w26 , w193 );
nor ( w195 , w194 , g3 );
nor ( w196 , w195 , w190 );
and ( w197 , w196 , w41 );
nor ( w198 , w197 , w176 );
not ( w199 , w15 );
and ( w200 , w199 , w198 );
not ( w201 , w25 );
and ( w202 , w200 , w201 );
or ( t_0 , w202 , w193 );

endmodule
