module patch (t_0, g1, g2);
input g1, g2;
output t_0;

or ( t_0 , g1 , g2 );

endmodule
