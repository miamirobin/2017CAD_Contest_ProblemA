module patch (t_0, g1);
input g1;
output t_0;

not ( t_0 , g1 );

endmodule
