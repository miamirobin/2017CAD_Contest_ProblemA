module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 ; 
output g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
n2450 ; 
wire t_0 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( n158 , g157 ); 
buf ( n159 , g158 ); 
buf ( n160 , g159 ); 
buf ( n161 , g160 ); 
buf ( n162 , g161 ); 
buf ( n163 , g162 ); 
buf ( n164 , g163 ); 
buf ( n165 , g164 ); 
buf ( n166 , g165 ); 
buf ( n167 , g166 ); 
buf ( n168 , g167 ); 
buf ( n169 , g168 ); 
buf ( n170 , g169 ); 
buf ( n171 , g170 ); 
buf ( n172 , g171 ); 
buf ( n173 , g172 ); 
buf ( n174 , g173 ); 
buf ( n175 , g174 ); 
buf ( n176 , g175 ); 
buf ( n177 , g176 ); 
buf ( n178 , g177 ); 
buf ( n179 , g178 ); 
buf ( g179 , n180 ); 
buf ( g180 , n181 ); 
buf ( g181 , n182 ); 
buf ( g182 , n183 ); 
buf ( g183 , n184 ); 
buf ( g184 , n185 ); 
buf ( g185 , n186 ); 
buf ( g186 , n187 ); 
buf ( g187 , n188 ); 
buf ( g188 , n189 ); 
buf ( g189 , n190 ); 
buf ( g190 , n191 ); 
buf ( g191 , n192 ); 
buf ( g192 , n193 ); 
buf ( g193 , n194 ); 
buf ( g194 , n195 ); 
buf ( g195 , n196 ); 
buf ( g196 , n197 ); 
buf ( g197 , n198 ); 
buf ( g198 , n199 ); 
buf ( g199 , n200 ); 
buf ( g200 , n201 ); 
buf ( g201 , n202 ); 
buf ( g202 , n203 ); 
buf ( g203 , n204 ); 
buf ( g204 , n205 ); 
buf ( g205 , n206 ); 
buf ( g206 , n207 ); 
buf ( g207 , n208 ); 
buf ( g208 , n209 ); 
buf ( g209 , n210 ); 
buf ( g210 , n211 ); 
buf ( g211 , n212 ); 
buf ( g212 , n213 ); 
buf ( g213 , n214 ); 
buf ( g214 , n215 ); 
buf ( g215 , n216 ); 
buf ( g216 , n217 ); 
buf ( g217 , n218 ); 
buf ( g218 , n219 ); 
buf ( g219 , n220 ); 
buf ( g220 , n221 ); 
buf ( g221 , n222 ); 
buf ( g222 , n223 ); 
buf ( g223 , n224 ); 
buf ( g224 , n225 ); 
buf ( g225 , n226 ); 
buf ( g226 , n227 ); 
buf ( g227 , n228 ); 
buf ( g228 , n229 ); 
buf ( g229 , n230 ); 
buf ( g230 , n231 ); 
buf ( g231 , n232 ); 
buf ( g232 , n233 ); 
buf ( g233 , n234 ); 
buf ( g234 , n235 ); 
buf ( g235 , n236 ); 
buf ( g236 , n237 ); 
buf ( g237 , n238 ); 
buf ( g238 , n239 ); 
buf ( g239 , n240 ); 
buf ( g240 , n241 ); 
buf ( g241 , n242 ); 
buf ( g242 , n243 ); 
buf ( n180 , n1807 ); 
buf ( n181 , n1999 ); 
buf ( n182 , n1851 ); 
buf ( n183 , n1452 ); 
buf ( n184 , n1795 ); 
buf ( n185 , n1508 ); 
buf ( n186 , n1989 ); 
buf ( n187 , n1266 ); 
buf ( n188 , n1559 ); 
buf ( n189 , n1337 ); 
buf ( n190 , n1691 ); 
buf ( n191 , n2450 ); 
buf ( n192 , n1858 ); 
buf ( n193 , n1567 ); 
buf ( n194 , n1606 ); 
buf ( n195 , n1615 ); 
buf ( n196 , n1896 ); 
buf ( n197 , n1343 ); 
buf ( n198 , n1786 ); 
buf ( n199 , n1347 ); 
buf ( n200 , n1695 ); 
buf ( n201 , n1770 ); 
buf ( n202 , n1901 ); 
buf ( n203 , n1700 ); 
buf ( n204 , n1705 ); 
buf ( n205 , n1710 ); 
buf ( n206 , n1963 ); 
buf ( n207 , n2352 ); 
buf ( n208 , n2306 ); 
buf ( n209 , n2392 ); 
buf ( n210 , n2397 ); 
buf ( n211 , n2440 ); 
buf ( n212 , n1980 ); 
buf ( n213 , n1944 ); 
buf ( n214 , n2060 ); 
buf ( n215 , n2022 ); 
buf ( n216 , n1924 ); 
buf ( n217 , n1781 ); 
buf ( n218 , n1916 ); 
buf ( n219 , n1653 ); 
buf ( n220 , n1958 ); 
buf ( n221 , n2153 ); 
buf ( n222 , n2326 ); 
buf ( n223 , n2367 ); 
buf ( n224 , n2313 ); 
buf ( n225 , n2372 ); 
buf ( n226 , n2404 ); 
buf ( n227 , n2331 ); 
buf ( n228 , n2436 ); 
buf ( n229 , n2141 ); 
buf ( n230 , n2257 ); 
buf ( n231 , n2217 ); 
buf ( n232 , n2147 ); 
buf ( n233 , n2346 ); 
buf ( n234 , n2385 ); 
buf ( n235 , n2266 ); 
buf ( n236 , n2389 ); 
buf ( n237 , n2445 ); 
buf ( n238 , n2095 ); 
buf ( n239 , n2198 ); 
buf ( n240 , n2301 ); 
buf ( n241 , n2427 ); 
buf ( n242 , n2432 ); 
buf ( n243 , n2425 ); 
nor ( n246 , n3 , n10 ); 
nor ( n247 , n9 , n23 ); 
nor ( n248 , n11 , n21 ); 
not ( n249 , n6 ); 
and ( n250 , n246 , n247 , n248 , n249 ); 
nor ( n251 , n2 , n5 ); 
nor ( n252 , n28 , n30 ); 
and ( n253 , n251 , n252 ); 
nand ( n254 , n250 , n253 ); 
and ( n255 , n1 , n24 , n26 ); 
and ( n256 , n254 , n255 ); 
nor ( n257 , n24 , n26 ); 
not ( n258 , n257 ); 
nor ( n259 , n258 , n1 ); 
nor ( n260 , n256 , n259 ); 
nor ( n261 , n2 , n23 , n28 ); 
nor ( n262 , n16 , n29 ); 
nand ( n263 , n261 , n262 , n257 ); 
nor ( n264 , n15 , n19 ); 
nor ( n265 , n6 , n21 ); 
nor ( n266 , n9 , n30 ); 
not ( n267 , n5 ); 
nand ( n268 , n264 , n265 , n266 , n267 ); 
nor ( n269 , n263 , n268 ); 
nor ( n270 , n18 , n20 ); 
nor ( n271 , n4 , n32 ); 
nor ( n272 , n12 , n22 ); 
not ( n273 , n11 ); 
nand ( n274 , n270 , n271 , n272 , n273 ); 
nor ( n275 , n3 , n13 ); 
nor ( n276 , n7 , n14 ); 
nor ( n277 , n10 , n17 ); 
nor ( n278 , n8 , n31 ); 
nand ( n279 , n275 , n276 , n277 , n278 ); 
nor ( n280 , n274 , n279 ); 
nand ( n281 , n269 , n280 ); 
nor ( n282 , n15 , n18 ); 
nor ( n283 , n19 , n20 ); 
nor ( n284 , n4 , n32 ); 
nand ( n285 , n282 , n283 , n262 , n284 ); 
nor ( n286 , n12 , n13 ); 
nor ( n287 , n14 , n17 ); 
nor ( n288 , n7 , n8 ); 
nor ( n289 , n22 , n31 ); 
nand ( n290 , n286 , n287 , n288 , n289 ); 
or ( n291 , n285 , n290 ); 
nand ( n292 , n291 , n255 ); 
nand ( n293 , n260 , n281 , n292 ); 
buf ( n294 , n293 ); 
not ( n295 , n294 ); 
not ( n296 , n168 ); 
and ( n297 , n295 , n296 ); 
not ( n298 , n295 ); 
not ( n299 , n3 ); 
not ( n300 , n299 ); 
not ( n301 , n2 ); 
not ( n302 , n301 ); 
not ( n303 , n9 ); 
nor ( n304 , n6 , n7 ); 
not ( n305 , n8 ); 
and ( n306 , n304 , n305 ); 
nand ( n307 , n303 , n306 ); 
nand ( n308 , n307 , n1 ); 
not ( n309 , n308 ); 
or ( n310 , n302 , n309 ); 
nand ( n311 , n310 , n1 ); 
not ( n312 , n311 ); 
or ( n313 , n300 , n312 ); 
or ( n314 , n311 , n299 ); 
nand ( n315 , n313 , n314 ); 
and ( n316 , n298 , n315 ); 
nor ( n317 , n297 , n316 ); 
xor ( n318 , n1 , n25 ); 
not ( n319 , n1 ); 
not ( n320 , n27 ); 
and ( n321 , n319 , n320 ); 
and ( n322 , n1 , n27 ); 
nor ( n323 , n321 , n322 ); 
nor ( n324 , n318 , n323 ); 
buf ( n325 , n324 ); 
and ( n326 , n325 , n52 ); 
not ( n327 , n323 ); 
and ( n328 , n1 , n25 ); 
nor ( n329 , n1 , n25 ); 
nor ( n330 , n328 , n329 ); 
nand ( n331 , n327 , n330 ); 
not ( n332 , n50 ); 
nor ( n333 , n331 , n332 ); 
nor ( n334 , n326 , n333 ); 
not ( n335 , n1 ); 
not ( n336 , n25 ); 
and ( n337 , n335 , n336 ); 
and ( n338 , n1 , n25 ); 
nor ( n339 , n337 , n338 ); 
not ( n340 , n339 ); 
xor ( n341 , n1 , n27 ); 
nand ( n342 , n340 , n341 ); 
not ( n343 , n342 ); 
and ( n344 , n343 , n49 ); 
not ( n345 , n51 ); 
xor ( n346 , n1 , n25 ); 
nand ( n347 , n346 , n341 ); 
buf ( n348 , n347 ); 
nor ( n349 , n345 , n348 ); 
nor ( n350 , n344 , n349 ); 
nand ( n351 , n334 , n350 ); 
buf ( n352 , n351 ); 
nor ( n353 , n317 , n352 ); 
not ( n354 , n353 ); 
nand ( n355 , n317 , n352 ); 
nand ( n356 , n354 , n355 ); 
not ( n357 , n356 ); 
buf ( n358 , n294 ); 
not ( n359 , n358 ); 
not ( n360 , n169 ); 
and ( n361 , n359 , n360 ); 
not ( n362 , n294 ); 
not ( n363 , n362 ); 
and ( n364 , n308 , n301 ); 
not ( n365 , n308 ); 
and ( n366 , n365 , n2 ); 
or ( n367 , n364 , n366 ); 
and ( n368 , n363 , n367 ); 
nor ( n369 , n361 , n368 ); 
and ( n370 , n325 , n45 ); 
not ( n371 , n46 ); 
xnor ( n372 , n1 , n27 ); 
nand ( n373 , n372 , n330 ); 
nor ( n374 , n371 , n373 ); 
nor ( n375 , n370 , n374 ); 
not ( n376 , n348 ); 
not ( n377 , n47 ); 
not ( n378 , n377 ); 
and ( n379 , n376 , n378 ); 
and ( n380 , n343 , n48 ); 
nor ( n381 , n379 , n380 ); 
nand ( n382 , n375 , n381 ); 
buf ( n383 , n382 ); 
not ( n384 , n383 ); 
or ( n385 , n369 , n384 ); 
nand ( n386 , n357 , n385 ); 
not ( n387 , n386 ); 
not ( n388 , n317 ); 
nand ( n389 , n352 , n388 ); 
not ( n390 , n389 ); 
not ( n391 , n342 ); 
and ( n392 , n391 , n33 ); 
not ( n393 , n331 ); 
and ( n394 , n393 , n34 ); 
nor ( n395 , n392 , n394 ); 
not ( n396 , n348 ); 
and ( n397 , n396 , n35 ); 
and ( n398 , n325 , n36 ); 
nor ( n399 , n397 , n398 ); 
nand ( n400 , n395 , n399 ); 
buf ( n401 , n400 ); 
nor ( n402 , n2 , n3 ); 
not ( n403 , n402 ); 
nand ( n404 , n403 , n1 ); 
nand ( n405 , n308 , n404 ); 
and ( n406 , n405 , n267 ); 
not ( n407 , n405 ); 
and ( n408 , n407 , n5 ); 
nor ( n409 , n406 , n408 ); 
not ( n410 , n409 ); 
not ( n411 , n358 ); 
or ( n412 , n410 , n411 ); 
not ( n413 , n171 ); 
nand ( n414 , n413 , n295 ); 
nand ( n415 , n412 , n414 ); 
xor ( n416 , n401 , n415 ); 
not ( n417 , n416 ); 
or ( n418 , n390 , n417 ); 
or ( n419 , n389 , n416 ); 
nand ( n420 , n418 , n419 ); 
not ( n421 , n420 ); 
or ( n422 , n387 , n421 ); 
not ( n423 , n416 ); 
or ( n424 , n423 , n389 ); 
nand ( n425 , n422 , n424 ); 
and ( n426 , n401 , n415 ); 
not ( n427 , n426 ); 
nor ( n428 , n358 , n166 ); 
not ( n429 , n428 ); 
buf ( n430 , n294 ); 
not ( n431 , n405 ); 
not ( n432 , n431 ); 
not ( n433 , n267 ); 
or ( n434 , n432 , n433 ); 
nand ( n435 , n434 , n1 ); 
not ( n436 , n4 ); 
nand ( n437 , n430 , n435 , n436 ); 
not ( n438 , n307 ); 
and ( n439 , n438 , n404 , n267 ); 
nand ( n440 , n1 , n4 ); 
nor ( n441 , n439 , n440 ); 
nand ( n442 , n363 , n441 ); 
nand ( n443 , n429 , n437 , n442 ); 
and ( n444 , n391 , n42 ); 
not ( n445 , n373 ); 
and ( n446 , n445 , n41 ); 
nor ( n447 , n444 , n446 ); 
not ( n448 , n348 ); 
not ( n449 , n43 ); 
not ( n450 , n449 ); 
and ( n451 , n448 , n450 ); 
and ( n452 , n325 , n44 ); 
nor ( n453 , n451 , n452 ); 
nand ( n454 , n447 , n453 ); 
buf ( n455 , n454 ); 
and ( n456 , n443 , n455 ); 
not ( n457 , n456 ); 
not ( n458 , n443 ); 
not ( n459 , n455 ); 
nand ( n460 , n458 , n459 ); 
nand ( n461 , n457 , n460 ); 
not ( n462 , n461 ); 
or ( n463 , n427 , n462 ); 
or ( n464 , n426 , n461 ); 
nand ( n465 , n463 , n464 ); 
and ( n466 , n425 , n465 ); 
not ( n467 , n426 ); 
nor ( n468 , n467 , n461 ); 
nor ( n469 , n466 , n468 ); 
and ( n470 , n251 , n299 , n436 ); 
nand ( n471 , n438 , n470 ); 
not ( n472 , n471 ); 
nor ( n473 , n472 , n273 ); 
not ( n474 , n473 ); 
nand ( n475 , n294 , n1 ); 
not ( n476 , n475 ); 
not ( n477 , n476 ); 
or ( n478 , n474 , n477 ); 
not ( n479 , n430 ); 
not ( n480 , n479 ); 
nor ( n481 , n471 , n11 ); 
and ( n482 , n480 , n481 ); 
not ( n483 , n165 ); 
not ( n484 , n483 ); 
not ( n485 , n295 ); 
or ( n486 , n484 , n485 ); 
not ( n487 , n1 ); 
nand ( n488 , n487 , n257 ); 
not ( n489 , n488 ); 
nand ( n490 , n489 , n273 ); 
nand ( n491 , n486 , n490 ); 
nor ( n492 , n482 , n491 ); 
nand ( n493 , n478 , n492 ); 
and ( n494 , n343 , n65 ); 
and ( n495 , n393 , n66 ); 
nor ( n496 , n494 , n495 ); 
not ( n497 , n347 ); 
and ( n498 , n497 , n67 ); 
and ( n499 , n325 , n68 ); 
nor ( n500 , n498 , n499 ); 
nand ( n501 , n496 , n500 ); 
buf ( n502 , n501 ); 
not ( n503 , n502 ); 
not ( n504 , n503 ); 
nand ( n505 , n493 , n504 ); 
not ( n506 , n505 ); 
not ( n507 , n10 ); 
or ( n508 , n481 , n507 ); 
nor ( n509 , n5 , n7 ); 
and ( n510 , n402 , n509 ); 
nor ( n511 , n4 , n8 ); 
nor ( n512 , n10 , n11 ); 
and ( n513 , n511 , n512 ); 
nor ( n514 , n6 , n9 ); 
nand ( n515 , n510 , n513 , n514 ); 
nand ( n516 , n508 , n515 ); 
not ( n517 , n516 ); 
not ( n518 , n476 ); 
or ( n519 , n517 , n518 ); 
nor ( n520 , n358 , n164 ); 
nor ( n521 , n488 , n10 ); 
nor ( n522 , n520 , n521 ); 
nand ( n523 , n519 , n522 ); 
buf ( n524 , n391 ); 
and ( n525 , n524 , n61 ); 
not ( n526 , n331 ); 
and ( n527 , n526 , n62 ); 
nor ( n528 , n525 , n527 ); 
not ( n529 , n348 ); 
and ( n530 , n529 , n63 ); 
and ( n531 , n325 , n64 ); 
nor ( n532 , n530 , n531 ); 
nand ( n533 , n528 , n532 ); 
nand ( n534 , n523 , n533 ); 
not ( n535 , n534 ); 
nor ( n536 , n523 , n533 ); 
nor ( n537 , n535 , n536 ); 
not ( n538 , n537 ); 
not ( n539 , n538 ); 
or ( n540 , n506 , n539 ); 
buf ( n541 , n456 ); 
not ( n542 , n541 ); 
not ( n543 , n493 ); 
or ( n544 , n543 , n502 ); 
nand ( n545 , n543 , n504 ); 
nand ( n546 , n544 , n545 ); 
not ( n547 , n546 ); 
nand ( n548 , n542 , n547 ); 
nand ( n549 , n540 , n548 ); 
nor ( n550 , n469 , n549 ); 
not ( n551 , n385 ); 
nand ( n552 , n356 , n551 ); 
nand ( n553 , n552 , n424 ); 
nor ( n554 , n468 , n553 ); 
xor ( n555 , n383 , n369 ); 
not ( n556 , n555 ); 
not ( n557 , n529 ); 
nand ( n558 , n325 , n40 ); 
and ( n559 , n341 , n37 ); 
and ( n560 , n339 , n38 ); 
nor ( n561 , n559 , n560 ); 
nand ( n562 , n557 , n558 , n561 ); 
not ( n563 , n562 ); 
and ( n564 , n262 , n288 , n287 , n264 ); 
nor ( n565 , n13 , n31 ); 
and ( n566 , n270 , n272 , n284 , n565 ); 
and ( n567 , n514 , n246 , n273 ); 
nand ( n568 , n564 , n566 , n567 , n253 ); 
nand ( n569 , n568 , n1 ); 
or ( n570 , n569 , n26 ); 
and ( n571 , n26 , n24 ); 
not ( n572 , n26 ); 
not ( n573 , n24 ); 
not ( n574 , n573 ); 
nor ( n575 , n21 , n23 ); 
not ( n576 , n575 ); 
or ( n577 , n574 , n576 ); 
nand ( n578 , n577 , n1 ); 
and ( n579 , n572 , n578 ); 
or ( n580 , n571 , n579 ); 
nand ( n581 , n570 , n580 ); 
not ( n582 , n575 ); 
and ( n583 , n582 , n1 ); 
nor ( n584 , n583 , n573 ); 
and ( n585 , n569 , n584 ); 
nor ( n586 , n581 , n585 ); 
or ( n587 , n170 , n586 ); 
not ( n588 , n9 ); 
or ( n589 , n306 , n487 , n588 ); 
not ( n590 , n308 ); 
or ( n591 , n590 , n9 ); 
nand ( n592 , n589 , n591 ); 
nand ( n593 , n586 , n592 ); 
nand ( n594 , n587 , n593 ); 
and ( n595 , n497 , n39 ); 
not ( n596 , n595 ); 
and ( n597 , n562 , n596 ); 
not ( n598 , n597 ); 
nor ( n599 , n594 , n598 ); 
nor ( n600 , n563 , n599 ); 
nand ( n601 , n556 , n600 ); 
not ( n602 , n601 ); 
and ( n603 , n343 , n155 ); 
and ( n604 , n325 , n156 ); 
nor ( n605 , n603 , n604 ); 
and ( n606 , n529 , n154 ); 
and ( n607 , n445 , n157 ); 
nor ( n608 , n606 , n607 ); 
nand ( n609 , n605 , n608 ); 
not ( n610 , n609 ); 
not ( n611 , n610 ); 
nor ( n612 , n487 , n304 ); 
xor ( n613 , n8 , n612 ); 
and ( n614 , n430 , n613 ); 
not ( n615 , n430 ); 
and ( n616 , n615 , n172 ); 
nor ( n617 , n614 , n616 ); 
nor ( n618 , n611 , n617 ); 
and ( n619 , n1 , n6 , n7 ); 
or ( n620 , n1 , n7 ); 
not ( n621 , n304 ); 
nand ( n622 , n620 , n621 ); 
nor ( n623 , n619 , n622 ); 
not ( n624 , n623 ); 
not ( n625 , n358 ); 
or ( n626 , n624 , n625 ); 
not ( n627 , n173 ); 
or ( n628 , n627 , n358 ); 
nand ( n629 , n626 , n628 ); 
and ( n630 , n391 , n153 ); 
and ( n631 , n445 , n152 ); 
nor ( n632 , n630 , n631 ); 
and ( n633 , n529 , n150 ); 
and ( n634 , n325 , n151 ); 
nor ( n635 , n633 , n634 ); 
nand ( n636 , n632 , n635 ); 
not ( n637 , n636 ); 
nand ( n638 , n629 , n637 ); 
not ( n639 , n638 ); 
nor ( n640 , n618 , n639 ); 
not ( n641 , n640 ); 
not ( n642 , n636 ); 
not ( n643 , n627 ); 
not ( n644 , n362 ); 
or ( n645 , n643 , n644 ); 
not ( n646 , n623 ); 
nand ( n647 , n646 , n358 ); 
nand ( n648 , n645 , n647 ); 
not ( n649 , n648 ); 
or ( n650 , n642 , n649 ); 
nand ( n651 , n650 , n638 ); 
not ( n652 , n651 ); 
not ( n653 , n249 ); 
not ( n654 , n358 ); 
or ( n655 , n653 , n654 ); 
not ( n656 , n174 ); 
nand ( n657 , n656 , n362 ); 
nand ( n658 , n655 , n657 ); 
not ( n659 , n147 ); 
not ( n660 , n391 ); 
or ( n661 , n659 , n660 ); 
nand ( n662 , n325 , n149 ); 
nand ( n663 , n661 , n662 ); 
not ( n664 , n146 ); 
not ( n665 , n497 ); 
or ( n666 , n664 , n665 ); 
nand ( n667 , n445 , n148 ); 
nand ( n668 , n666 , n667 ); 
nor ( n669 , n663 , n668 ); 
not ( n670 , n669 ); 
nor ( n671 , n658 , n670 ); 
nand ( n672 , n652 , n671 ); 
not ( n673 , n672 ); 
or ( n674 , n641 , n673 ); 
not ( n675 , n617 ); 
not ( n676 , n675 ); 
nand ( n677 , n676 , n611 ); 
nand ( n678 , n674 , n677 ); 
not ( n679 , n678 ); 
not ( n680 , n679 ); 
or ( n681 , n602 , n680 ); 
and ( n682 , n594 , n597 ); 
not ( n683 , n594 ); 
and ( n684 , n683 , n598 ); 
nor ( n685 , n682 , n684 ); 
not ( n686 , n685 ); 
and ( n687 , n601 , n686 ); 
nor ( n688 , n556 , n600 ); 
nor ( n689 , n687 , n688 ); 
nand ( n690 , n681 , n689 ); 
nand ( n691 , n554 , n690 ); 
and ( n692 , n524 , n53 ); 
buf ( n693 , n325 ); 
and ( n694 , n693 , n56 ); 
nor ( n695 , n692 , n694 ); 
not ( n696 , n557 ); 
not ( n697 , n55 ); 
not ( n698 , n697 ); 
and ( n699 , n696 , n698 ); 
and ( n700 , n526 , n54 ); 
nor ( n701 , n699 , n700 ); 
nand ( n702 , n695 , n701 ); 
nor ( n703 , n515 , n13 ); 
not ( n704 , n12 ); 
or ( n705 , n703 , n704 ); 
and ( n706 , n514 , n286 ); 
nand ( n707 , n706 , n510 , n513 ); 
buf ( n708 , n707 ); 
nand ( n709 , n705 , n708 ); 
not ( n710 , n709 ); 
not ( n711 , n476 ); 
or ( n712 , n710 , n711 ); 
not ( n713 , n363 ); 
not ( n714 , n163 ); 
and ( n715 , n713 , n714 ); 
nor ( n716 , n488 , n12 ); 
nor ( n717 , n715 , n716 ); 
nand ( n718 , n712 , n717 ); 
nand ( n719 , n702 , n718 ); 
not ( n720 , n14 ); 
not ( n721 , n708 ); 
or ( n722 , n720 , n721 ); 
or ( n723 , n708 , n14 ); 
nand ( n724 , n722 , n723 ); 
not ( n725 , n724 ); 
not ( n726 , n476 ); 
or ( n727 , n725 , n726 ); 
nor ( n728 , n358 , n162 ); 
nor ( n729 , n488 , n14 ); 
nor ( n730 , n728 , n729 ); 
nand ( n731 , n727 , n730 ); 
and ( n732 , n524 , n69 ); 
and ( n733 , n526 , n70 ); 
nor ( n734 , n732 , n733 ); 
and ( n735 , n529 , n71 ); 
and ( n736 , n693 , n72 ); 
nor ( n737 , n735 , n736 ); 
nand ( n738 , n734 , n737 ); 
nor ( n739 , n731 , n738 ); 
not ( n740 , n739 ); 
nand ( n741 , n731 , n738 ); 
nand ( n742 , n740 , n741 ); 
nand ( n743 , n719 , n742 ); 
not ( n744 , n16 ); 
not ( n745 , n723 ); 
or ( n746 , n744 , n745 ); 
or ( n747 , n14 , n16 ); 
nor ( n748 , n707 , n747 ); 
not ( n749 , n748 ); 
nand ( n750 , n746 , n749 ); 
not ( n751 , n750 ); 
not ( n752 , n476 ); 
or ( n753 , n751 , n752 ); 
nor ( n754 , n363 , n177 ); 
nor ( n755 , n488 , n16 ); 
nor ( n756 , n754 , n755 ); 
nand ( n757 , n753 , n756 ); 
and ( n758 , n524 , n73 ); 
and ( n759 , n693 , n76 ); 
nor ( n760 , n758 , n759 ); 
and ( n761 , n529 , n75 ); 
and ( n762 , n526 , n74 ); 
nor ( n763 , n761 , n762 ); 
nand ( n764 , n760 , n763 ); 
or ( n765 , n757 , n764 ); 
nand ( n766 , n757 , n764 ); 
nand ( n767 , n765 , n766 ); 
nand ( n768 , n767 , n741 ); 
and ( n769 , n743 , n768 ); 
not ( n770 , n718 ); 
not ( n771 , n702 ); 
not ( n772 , n771 ); 
or ( n773 , n770 , n772 ); 
not ( n774 , n718 ); 
nand ( n775 , n774 , n702 ); 
nand ( n776 , n773 , n775 ); 
not ( n777 , n776 ); 
and ( n778 , n515 , n13 ); 
nor ( n779 , n778 , n703 ); 
not ( n780 , n779 ); 
not ( n781 , n780 ); 
not ( n782 , n476 ); 
or ( n783 , n781 , n782 ); 
not ( n784 , n488 ); 
not ( n785 , n13 ); 
and ( n786 , n784 , n785 ); 
not ( n787 , n167 ); 
and ( n788 , n479 , n787 ); 
nor ( n789 , n786 , n788 ); 
nand ( n790 , n783 , n789 ); 
and ( n791 , n524 , n58 ); 
and ( n792 , n526 , n59 ); 
nor ( n793 , n791 , n792 ); 
and ( n794 , n529 , n57 ); 
and ( n795 , n325 , n60 ); 
nor ( n796 , n794 , n795 ); 
nand ( n797 , n793 , n796 ); 
nand ( n798 , n790 , n797 ); 
nand ( n799 , n777 , n798 ); 
nor ( n800 , n790 , n797 ); 
not ( n801 , n800 ); 
nand ( n802 , n801 , n798 ); 
buf ( n803 , n534 ); 
nand ( n804 , n802 , n803 ); 
not ( n805 , n17 ); 
not ( n806 , n749 ); 
or ( n807 , n805 , n806 ); 
not ( n808 , n17 ); 
nand ( n809 , n808 , n748 ); 
nand ( n810 , n807 , n809 ); 
not ( n811 , n810 ); 
not ( n812 , n476 ); 
or ( n813 , n811 , n812 ); 
not ( n814 , n295 ); 
nor ( n815 , n814 , n176 ); 
nor ( n816 , n488 , n17 ); 
nor ( n817 , n815 , n816 ); 
nand ( n818 , n813 , n817 ); 
not ( n819 , n818 ); 
not ( n820 , n819 ); 
and ( n821 , n529 , n83 ); 
and ( n822 , n524 , n81 ); 
nor ( n823 , n821 , n822 ); 
buf ( n824 , n526 ); 
and ( n825 , n824 , n82 ); 
and ( n826 , n693 , n84 ); 
nor ( n827 , n825 , n826 ); 
nand ( n828 , n823 , n827 ); 
not ( n829 , n828 ); 
and ( n830 , n820 , n829 ); 
not ( n831 , n828 ); 
nor ( n832 , n831 , n818 ); 
nor ( n833 , n830 , n832 ); 
nand ( n834 , n833 , n766 ); 
and ( n835 , n769 , n799 , n804 , n834 ); 
nand ( n836 , n550 , n691 , n835 ); 
not ( n837 , n766 ); 
buf ( n838 , n833 ); 
not ( n839 , n838 ); 
nand ( n840 , n837 , n839 ); 
nand ( n841 , n836 , n840 ); 
nand ( n842 , n818 , n828 ); 
and ( n843 , n841 , n842 ); 
not ( n844 , n841 ); 
not ( n845 , n536 ); 
not ( n846 , n845 ); 
not ( n847 , n503 ); 
not ( n848 , n543 ); 
or ( n849 , n847 , n848 ); 
nand ( n850 , n849 , n541 ); 
nand ( n851 , n850 , n505 ); 
not ( n852 , n851 ); 
or ( n853 , n846 , n852 ); 
nand ( n854 , n853 , n803 ); 
not ( n855 , n802 ); 
nand ( n856 , n854 , n855 ); 
not ( n857 , n856 ); 
not ( n858 , n719 ); 
not ( n859 , n742 ); 
nand ( n860 , n858 , n859 ); 
buf ( n861 , n741 ); 
and ( n862 , n860 , n861 , n798 ); 
not ( n863 , n862 ); 
or ( n864 , n857 , n863 ); 
not ( n865 , n719 ); 
not ( n866 , n777 ); 
or ( n867 , n865 , n866 ); 
not ( n868 , n739 ); 
nand ( n869 , n867 , n868 ); 
and ( n870 , n869 , n861 ); 
not ( n871 , n767 ); 
not ( n872 , n871 ); 
nor ( n873 , n870 , n872 ); 
nand ( n874 , n864 , n873 ); 
and ( n875 , n874 , n842 ); 
and ( n876 , n819 , n831 ); 
nor ( n877 , n875 , n876 ); 
and ( n878 , n844 , n877 ); 
nor ( n879 , n843 , n878 ); 
not ( n880 , n28 ); 
not ( n881 , n880 ); 
not ( n882 , n29 ); 
not ( n883 , n32 ); 
and ( n884 , n264 , n270 , n808 ); 
nand ( n885 , n882 , n883 , n748 , n884 ); 
not ( n886 , n885 ); 
not ( n887 , n886 ); 
or ( n888 , n881 , n887 ); 
nand ( n889 , n888 , n30 ); 
not ( n890 , n889 ); 
buf ( n891 , n252 ); 
and ( n892 , n886 , n891 ); 
nor ( n893 , n892 , n487 ); 
not ( n894 , n893 ); 
or ( n895 , n890 , n894 ); 
nand ( n896 , n487 , n30 ); 
nand ( n897 , n895 , n896 ); 
and ( n898 , n748 , n884 ); 
nand ( n899 , n1 , n29 ); 
or ( n900 , n898 , n899 ); 
or ( n901 , n1 , n29 ); 
nand ( n902 , n900 , n901 ); 
not ( n903 , n29 ); 
and ( n904 , n748 , n884 , n903 ); 
or ( n905 , n902 , n904 ); 
and ( n906 , n897 , n905 ); 
not ( n907 , n897 ); 
not ( n908 , n32 ); 
nor ( n909 , n904 , n908 ); 
nand ( n910 , n885 , n1 ); 
or ( n911 , n909 , n910 ); 
or ( n912 , n908 , n1 ); 
nand ( n913 , n911 , n912 ); 
not ( n914 , n913 ); 
and ( n915 , n907 , n914 ); 
nor ( n916 , n906 , n915 ); 
not ( n917 , n916 ); 
not ( n918 , n28 ); 
not ( n919 , n910 ); 
or ( n920 , n918 , n919 ); 
or ( n921 , n910 , n28 ); 
nand ( n922 , n920 , n921 ); 
and ( n923 , n897 , n922 ); 
not ( n924 , n923 ); 
not ( n925 , n897 ); 
not ( n926 , n922 ); 
nand ( n927 , n925 , n926 ); 
nand ( n928 , n924 , n927 ); 
nor ( n929 , n917 , n928 ); 
not ( n930 , n929 ); 
not ( n931 , n930 ); 
buf ( n932 , n931 ); 
not ( n933 , n932 ); 
and ( n934 , n524 , n78 ); 
and ( n935 , n693 , n80 ); 
nor ( n936 , n934 , n935 ); 
and ( n937 , n529 , n77 ); 
and ( n938 , n824 , n79 ); 
nor ( n939 , n937 , n938 ); 
nand ( n940 , n936 , n939 ); 
not ( n941 , n480 ); 
not ( n942 , n175 ); 
and ( n943 , n941 , n942 ); 
not ( n944 , n809 ); 
nand ( n945 , n944 , n480 ); 
and ( n946 , n945 , n488 ); 
nor ( n947 , n946 , n15 ); 
nor ( n948 , n943 , n947 ); 
nand ( n949 , n476 , n809 , n15 ); 
and ( n950 , n948 , n949 ); 
and ( n951 , n940 , n950 ); 
not ( n952 , n940 ); 
not ( n953 , n950 ); 
and ( n954 , n952 , n953 ); 
nor ( n955 , n951 , n954 ); 
buf ( n956 , n955 ); 
nor ( n957 , n933 , n956 ); 
and ( n958 , n879 , n957 ); 
not ( n959 , n879 ); 
and ( n960 , n932 , n956 ); 
and ( n961 , n959 , n960 ); 
nor ( n962 , n958 , n961 ); 
nor ( n963 , n928 , n916 ); 
buf ( n964 , n963 ); 
nand ( n965 , n964 , n955 ); 
not ( n966 , n965 ); 
not ( n967 , n742 ); 
nand ( n968 , n967 , n775 ); 
not ( n969 , n738 ); 
nor ( n970 , n731 , n969 ); 
not ( n971 , n970 ); 
nand ( n972 , n971 , n871 ); 
nand ( n973 , n968 , n972 ); 
not ( n974 , n523 ); 
and ( n975 , n974 , n533 ); 
not ( n976 , n975 ); 
not ( n977 , n976 ); 
not ( n978 , n855 ); 
or ( n979 , n977 , n978 ); 
not ( n980 , n790 ); 
nand ( n981 , n980 , n797 ); 
nand ( n982 , n776 , n981 ); 
nand ( n983 , n979 , n982 ); 
nor ( n984 , n973 , n983 ); 
not ( n985 , n984 ); 
nor ( n986 , n669 , n658 ); 
nor ( n987 , n986 , n636 ); 
nand ( n988 , n675 , n611 ); 
and ( n989 , n987 , n988 ); 
not ( n990 , n599 ); 
nand ( n991 , n598 , n594 ); 
nand ( n992 , n990 , n991 ); 
nor ( n993 , n989 , n992 ); 
not ( n994 , n610 ); 
not ( n995 , n617 ); 
or ( n996 , n994 , n995 ); 
nand ( n997 , n648 , n637 ); 
nand ( n998 , n996 , n997 ); 
not ( n999 , n670 ); 
and ( n1000 , n295 , n174 ); 
not ( n1001 , n295 ); 
and ( n1002 , n1001 , n6 ); 
nor ( n1003 , n1000 , n1002 ); 
nor ( n1004 , n999 , n1003 ); 
nor ( n1005 , n629 , n1004 ); 
or ( n1006 , n998 , n1005 ); 
nand ( n1007 , n1006 , n988 ); 
nand ( n1008 , n993 , n1007 ); 
buf ( n1009 , n595 ); 
nor ( n1010 , n1009 , n599 ); 
or ( n1011 , n556 , n1010 ); 
nand ( n1012 , n1008 , n1011 ); 
and ( n1013 , n383 , n369 ); 
xor ( n1014 , n356 , n1013 ); 
and ( n1015 , n556 , n1010 ); 
nor ( n1016 , n1014 , n1015 ); 
nand ( n1017 , n1012 , n1016 ); 
not ( n1018 , n1017 ); 
not ( n1019 , n415 ); 
and ( n1020 , n1019 , n401 ); 
nand ( n1021 , n461 , n1020 ); 
not ( n1022 , n1021 ); 
not ( n1023 , n355 ); 
nand ( n1024 , n1023 , n423 ); 
nand ( n1025 , n357 , n1013 ); 
nand ( n1026 , n1024 , n1025 ); 
nor ( n1027 , n1022 , n1026 ); 
not ( n1028 , n1027 ); 
or ( n1029 , n1018 , n1028 ); 
xor ( n1030 , n455 , n458 ); 
xor ( n1031 , n1030 , n1020 ); 
nand ( n1032 , n416 , n355 ); 
nand ( n1033 , n1031 , n1032 ); 
and ( n1034 , n1033 , n1021 ); 
and ( n1035 , n458 , n455 ); 
not ( n1036 , n1035 ); 
and ( n1037 , n546 , n1036 ); 
nor ( n1038 , n1034 , n1037 ); 
nand ( n1039 , n1029 , n1038 ); 
buf ( n1040 , n545 ); 
and ( n1041 , n537 , n1040 ); 
nor ( n1042 , n1039 , n1041 ); 
not ( n1043 , n1042 ); 
or ( n1044 , n985 , n1043 ); 
nand ( n1045 , n1044 , n839 ); 
not ( n1046 , n757 ); 
and ( n1047 , n1046 , n764 ); 
nand ( n1048 , n1045 , n1047 ); 
and ( n1049 , n1048 , n832 ); 
not ( n1050 , n1048 ); 
not ( n1051 , n832 ); 
and ( n1052 , n1050 , n1051 ); 
nor ( n1053 , n1049 , n1052 ); 
nand ( n1054 , n802 , n975 ); 
nand ( n1055 , n1041 , n1054 ); 
and ( n1056 , n984 , n1055 ); 
not ( n1057 , n1056 ); 
not ( n1058 , n1040 ); 
nand ( n1059 , n547 , n1035 ); 
not ( n1060 , n1059 ); 
or ( n1061 , n1058 , n1060 ); 
nand ( n1062 , n1061 , n538 ); 
and ( n1063 , n1062 , n1054 ); 
nand ( n1064 , n1039 , n1063 ); 
not ( n1065 , n1064 ); 
or ( n1066 , n1057 , n1065 ); 
not ( n1067 , n973 ); 
not ( n1068 , n981 ); 
nand ( n1069 , n1068 , n777 ); 
not ( n1070 , n1069 ); 
and ( n1071 , n1067 , n1070 ); 
or ( n1072 , n859 , n775 ); 
not ( n1073 , n872 ); 
or ( n1074 , n1072 , n1073 ); 
nand ( n1075 , n872 , n970 ); 
nand ( n1076 , n1074 , n1075 ); 
nor ( n1077 , n1071 , n1076 ); 
nand ( n1078 , n1066 , n1077 ); 
nand ( n1079 , n1078 , n838 ); 
nand ( n1080 , n966 , n1053 , n1079 ); 
buf ( n1081 , n569 ); 
buf ( n1082 , n1081 ); 
nand ( n1083 , n1082 , n578 ); 
not ( n1084 , n26 ); 
and ( n1085 , n1083 , n1084 ); 
not ( n1086 , n1083 ); 
and ( n1087 , n1086 , n26 ); 
or ( n1088 , n1085 , n1087 ); 
nand ( n1089 , n351 , n501 , n595 ); 
not ( n1090 , n1089 ); 
nand ( n1091 , n382 , n454 , n400 ); 
not ( n1092 , n1091 ); 
nand ( n1093 , n1090 , n1092 , n533 ); 
not ( n1094 , n1093 ); 
nand ( n1095 , n1094 , n797 , n702 ); 
nor ( n1096 , n1095 , n969 ); 
and ( n1097 , n1096 , n764 ); 
not ( n1098 , n1097 ); 
and ( n1099 , n1098 , n828 ); 
not ( n1100 , n1098 ); 
and ( n1101 , n1100 , n831 ); 
nor ( n1102 , n1099 , n1101 ); 
and ( n1103 , n1088 , n1102 ); 
not ( n1104 , n1088 ); 
nor ( n1105 , n1091 , n1089 ); 
or ( n1106 , n1105 , n533 ); 
nand ( n1107 , n1106 , n1093 ); 
not ( n1108 , n1107 ); 
and ( n1109 , n693 , n144 ); 
not ( n1110 , n145 ); 
not ( n1111 , n343 ); 
or ( n1112 , n1110 , n1111 ); 
nand ( n1113 , n445 , n143 ); 
nand ( n1114 , n1112 , n1113 ); 
nor ( n1115 , n1109 , n1114 ); 
nor ( n1116 , n669 , n1115 ); 
and ( n1117 , n1116 , n636 ); 
and ( n1118 , n597 , n609 ); 
nand ( n1119 , n1117 , n1118 ); 
nand ( n1120 , n401 , n502 , n383 , n352 ); 
nor ( n1121 , n1119 , n1120 ); 
not ( n1122 , n455 ); 
not ( n1123 , n351 ); 
nand ( n1124 , n382 , n595 ); 
nor ( n1125 , n1123 , n1124 ); 
nand ( n1126 , n1125 , n401 ); 
nand ( n1127 , n1122 , n1126 ); 
nand ( n1128 , n1108 , n1121 , n1127 ); 
nand ( n1129 , n702 , n797 ); 
nor ( n1130 , n1128 , n1129 ); 
nand ( n1131 , n1130 , n738 ); 
not ( n1132 , n1131 ); 
xnor ( n1133 , n1095 , n764 ); 
nand ( n1134 , n1132 , n1133 ); 
not ( n1135 , n1134 ); 
and ( n1136 , n940 , n828 ); 
nand ( n1137 , n1135 , n1136 ); 
nand ( n1138 , n1097 , n1136 ); 
and ( n1139 , n524 , n121 ); 
and ( n1140 , n824 , n122 ); 
nor ( n1141 , n1139 , n1140 ); 
and ( n1142 , n529 , n123 ); 
and ( n1143 , n693 , n120 ); 
nor ( n1144 , n1142 , n1143 ); 
nand ( n1145 , n1141 , n1144 ); 
not ( n1146 , n1145 ); 
and ( n1147 , n1138 , n1146 ); 
not ( n1148 , n1138 ); 
and ( n1149 , n1148 , n1145 ); 
nor ( n1150 , n1147 , n1149 ); 
xor ( n1151 , n1137 , n1150 ); 
and ( n1152 , n1104 , n1151 ); 
nor ( n1153 , n1103 , n1152 ); 
not ( n1154 , n923 ); 
buf ( n1155 , n1154 ); 
not ( n1156 , n1155 ); 
nand ( n1157 , n1153 , n1156 ); 
buf ( n1158 , n731 ); 
and ( n1159 , n1158 , n757 ); 
not ( n1160 , n980 ); 
not ( n1161 , n774 ); 
nand ( n1162 , n1159 , n1160 , n1161 , n818 ); 
not ( n1163 , n1162 ); 
not ( n1164 , n369 ); 
nand ( n1165 , n388 , n1164 ); 
not ( n1166 , n1165 ); 
not ( n1167 , n675 ); 
not ( n1168 , n1019 ); 
nand ( n1169 , n1167 , n1168 ); 
nand ( n1170 , n658 , n648 ); 
nor ( n1171 , n1169 , n1170 ); 
buf ( n1172 , n594 ); 
nand ( n1173 , n1166 , n1171 , n1172 ); 
not ( n1174 , n1173 ); 
nor ( n1175 , n543 , n458 ); 
nand ( n1176 , n1174 , n1175 ); 
nor ( n1177 , n1176 , n974 ); 
buf ( n1178 , n1177 ); 
nand ( n1179 , n1163 , n1178 ); 
and ( n1180 , n1179 , n950 ); 
not ( n1181 , n1179 ); 
and ( n1182 , n1181 , n953 ); 
nor ( n1183 , n1180 , n1182 ); 
not ( n1184 , n927 ); 
not ( n1185 , n913 ); 
nand ( n1186 , n1185 , n905 ); 
not ( n1187 , n1186 ); 
nand ( n1188 , n1184 , n1187 ); 
not ( n1189 , n1188 ); 
nand ( n1190 , n1183 , n1189 ); 
nand ( n1191 , n1184 , n913 ); 
not ( n1192 , n1191 ); 
nand ( n1193 , n1192 , n950 ); 
and ( n1194 , n1157 , n1190 , n1193 ); 
nand ( n1195 , n962 , n1080 , n1194 ); 
nand ( n1196 , n1053 , n1079 ); 
or ( n1197 , n928 , n916 ); 
buf ( n1198 , n1197 ); 
nor ( n1199 , n1198 , n956 ); 
nand ( n1200 , n1196 , n1199 ); 
not ( n1201 , n1200 ); 
nor ( n1202 , n1195 , n1201 ); 
not ( n1203 , n21 ); 
not ( n1204 , n1 ); 
or ( n1205 , n1203 , n1204 ); 
nand ( n1206 , n1205 , n1081 ); 
nand ( n1207 , n568 , n21 ); 
and ( n1208 , n1206 , n1207 ); 
and ( n1209 , n487 , n21 ); 
nor ( n1210 , n1208 , n1209 ); 
not ( n1211 , n1210 ); 
not ( n1212 , n31 ); 
not ( n1213 , n1212 ); 
not ( n1214 , n891 ); 
nor ( n1215 , n1214 , n885 ); 
not ( n1216 , n1215 ); 
or ( n1217 , n1213 , n1216 ); 
nand ( n1218 , n1217 , n22 ); 
not ( n1219 , n1082 ); 
and ( n1220 , n1218 , n1219 ); 
and ( n1221 , n487 , n22 ); 
nor ( n1222 , n1220 , n1221 ); 
not ( n1223 , n1222 ); 
xor ( n1224 , n1206 , n23 ); 
and ( n1225 , n1223 , n1224 ); 
nand ( n1226 , n1211 , n1225 ); 
xnor ( n1227 , n893 , n1212 ); 
not ( n1228 , n158 ); 
nor ( n1229 , n1227 , n1228 ); 
and ( n1230 , n1226 , n1229 ); 
nor ( n1231 , n1224 , n1210 ); 
not ( n1232 , n1231 ); 
not ( n1233 , n159 ); 
nand ( n1234 , n1225 , n1233 ); 
and ( n1235 , n1210 , n159 ); 
not ( n1236 , n1235 ); 
not ( n1237 , n1222 ); 
or ( n1238 , n1236 , n1237 ); 
not ( n1239 , n161 ); 
nand ( n1240 , n1238 , n1239 ); 
nand ( n1241 , n1240 , n1224 ); 
nand ( n1242 , n1232 , n1234 , n1241 ); 
not ( n1243 , n1242 ); 
not ( n1244 , n926 ); 
not ( n1245 , n925 ); 
not ( n1246 , n1245 ); 
or ( n1247 , n1244 , n1246 ); 
nand ( n1248 , n1247 , n1186 ); 
and ( n1249 , n926 , n914 ); 
nor ( n1250 , n1249 , n1245 ); 
nor ( n1251 , n1248 , n1250 ); 
not ( n1252 , n1251 ); 
nor ( n1253 , n1233 , n160 ); 
nand ( n1254 , n1225 , n1253 ); 
or ( n1255 , n1235 , n160 ); 
nand ( n1256 , n1255 , n1224 ); 
nand ( n1257 , n1256 , n1222 ); 
and ( n1258 , n1254 , n1257 ); 
not ( n1259 , n1258 ); 
and ( n1260 , n1230 , n1243 , n1252 , n1259 ); 
buf ( n1261 , n1260 ); 
not ( n1262 , n1261 ); 
or ( n1263 , n1202 , n1262 ); 
not ( n1264 , n80 ); 
or ( n1265 , n1261 , n1264 ); 
nand ( n1266 , n1263 , n1265 ); 
not ( n1267 , n1072 ); 
and ( n1268 , n1041 , n1054 ); 
nor ( n1269 , n1268 , n983 ); 
not ( n1270 , n1269 ); 
not ( n1271 , n1064 ); 
or ( n1272 , n1270 , n1271 ); 
nand ( n1273 , n1272 , n1069 ); 
nand ( n1274 , n1273 , n968 ); 
not ( n1275 , n1274 ); 
or ( n1276 , n1267 , n1275 ); 
and ( n1277 , n1075 , n972 ); 
nor ( n1278 , n1198 , n1277 ); 
nand ( n1279 , n1276 , n1278 ); 
and ( n1280 , n964 , n1277 , n1072 ); 
nand ( n1281 , n1274 , n1280 ); 
nand ( n1282 , n1279 , n1281 ); 
not ( n1283 , n1189 ); 
and ( n1284 , n1177 , n790 ); 
and ( n1285 , n1284 , n1161 ); 
and ( n1286 , n1285 , n1158 ); 
and ( n1287 , n1286 , n1046 ); 
not ( n1288 , n1286 ); 
not ( n1289 , n1046 ); 
and ( n1290 , n1288 , n1289 ); 
nor ( n1291 , n1287 , n1290 ); 
nor ( n1292 , n1283 , n1291 ); 
nor ( n1293 , n1282 , n1292 ); 
not ( n1294 , n1293 ); 
not ( n1295 , n932 ); 
and ( n1296 , n861 , n872 ); 
not ( n1297 , n861 ); 
and ( n1298 , n1297 , n1073 ); 
or ( n1299 , n1296 , n1298 ); 
buf ( n1300 , n860 ); 
not ( n1301 , n1300 ); 
and ( n1302 , n856 , n798 ); 
nor ( n1303 , n1302 , n777 ); 
nor ( n1304 , n1301 , n1303 ); 
not ( n1305 , n1304 ); 
and ( n1306 , n799 , n804 ); 
nand ( n1307 , n550 , n691 , n1306 ); 
not ( n1308 , n1307 ); 
or ( n1309 , n1305 , n1308 ); 
buf ( n1310 , n743 ); 
nand ( n1311 , n1309 , n1310 ); 
xor ( n1312 , n1299 , n1311 ); 
not ( n1313 , n1312 ); 
or ( n1314 , n1295 , n1313 ); 
not ( n1315 , n1135 ); 
not ( n1316 , n1315 ); 
not ( n1317 , n1102 ); 
or ( n1318 , n1316 , n1317 ); 
or ( n1319 , n831 , n1315 ); 
nand ( n1320 , n1318 , n1319 ); 
not ( n1321 , n1088 ); 
and ( n1322 , n1320 , n1321 ); 
not ( n1323 , n1088 ); 
buf ( n1324 , n1095 ); 
and ( n1325 , n1324 , n969 ); 
nor ( n1326 , n1325 , n1096 ); 
nor ( n1327 , n1323 , n1326 ); 
nor ( n1328 , n1322 , n1327 ); 
and ( n1329 , n1328 , n1156 ); 
and ( n1330 , n1192 , n1046 ); 
nor ( n1331 , n1329 , n1330 ); 
nand ( n1332 , n1314 , n1331 ); 
nor ( n1333 , n1294 , n1332 ); 
or ( n1334 , n1333 , n1262 ); 
not ( n1335 , n76 ); 
or ( n1336 , n1261 , n1335 ); 
nand ( n1337 , n1334 , n1336 ); 
and ( n1338 , n1230 , n1243 , n1258 , n1252 ); 
not ( n1339 , n1338 ); 
or ( n1340 , n1202 , n1339 ); 
not ( n1341 , n79 ); 
or ( n1342 , n1341 , n1338 ); 
nand ( n1343 , n1340 , n1342 ); 
or ( n1344 , n1333 , n1339 ); 
not ( n1345 , n74 ); 
or ( n1346 , n1345 , n1338 ); 
nand ( n1347 , n1344 , n1346 ); 
buf ( n1348 , n1031 ); 
not ( n1349 , n1348 ); 
not ( n1350 , n1025 ); 
not ( n1351 , n1017 ); 
or ( n1352 , n1350 , n1351 ); 
and ( n1353 , n1032 , n1024 ); 
nand ( n1354 , n1352 , n1353 ); 
nand ( n1355 , n1354 , n1024 ); 
not ( n1356 , n1355 ); 
or ( n1357 , n1349 , n1356 ); 
buf ( n1358 , n1021 ); 
nand ( n1359 , n1357 , n1358 ); 
not ( n1360 , n1359 ); 
buf ( n1361 , n1059 ); 
nand ( n1362 , n1360 , n1361 ); 
not ( n1363 , n1037 ); 
not ( n1364 , n1363 ); 
not ( n1365 , n538 ); 
and ( n1366 , n1040 , n1365 ); 
not ( n1367 , n1040 ); 
and ( n1368 , n1367 , n538 ); 
nor ( n1369 , n1366 , n1368 ); 
nor ( n1370 , n1197 , n1364 , n1369 ); 
and ( n1371 , n1362 , n1370 ); 
and ( n1372 , n505 , n1365 ); 
not ( n1373 , n505 ); 
and ( n1374 , n1373 , n538 ); 
nor ( n1375 , n1372 , n1374 ); 
not ( n1376 , n547 ); 
nand ( n1377 , n1376 , n541 ); 
not ( n1378 , n1377 ); 
not ( n1379 , n1378 ); 
not ( n1380 , n469 ); 
nand ( n1381 , n691 , n1380 , n548 ); 
nand ( n1382 , n1379 , n1381 ); 
xor ( n1383 , n1375 , n1382 ); 
nor ( n1384 , n1383 , n933 ); 
nor ( n1385 , n1371 , n1384 ); 
not ( n1386 , n1364 ); 
not ( n1387 , n1359 ); 
nand ( n1388 , n1387 , n1361 ); 
nand ( n1389 , n1386 , n1388 ); 
nand ( n1390 , n1389 , n964 , n1369 ); 
nand ( n1391 , n1385 , n1390 ); 
not ( n1392 , n1154 ); 
nand ( n1393 , n1392 , n1321 ); 
not ( n1394 , n1393 ); 
not ( n1395 , n1093 ); 
xor ( n1396 , n797 , n1395 ); 
not ( n1397 , n1396 ); 
buf ( n1398 , n1128 ); 
not ( n1399 , n1398 ); 
or ( n1400 , n1397 , n1399 ); 
or ( n1401 , n1398 , n797 ); 
nand ( n1402 , n1400 , n1401 ); 
and ( n1403 , n1394 , n1402 ); 
and ( n1404 , n923 , n1088 ); 
not ( n1405 , n1126 ); 
nand ( n1406 , n1405 , n455 ); 
and ( n1407 , n1406 , n503 ); 
not ( n1408 , n1406 ); 
and ( n1409 , n1408 , n504 ); 
nor ( n1410 , n1407 , n1409 ); 
and ( n1411 , n1404 , n1410 ); 
nor ( n1412 , n1403 , n1411 ); 
or ( n1413 , n1412 , n1186 ); 
not ( n1414 , n1178 ); 
and ( n1415 , n1176 , n974 ); 
not ( n1416 , n1189 ); 
nor ( n1417 , n1415 , n1416 ); 
nand ( n1418 , n1414 , n1417 ); 
nand ( n1419 , n1413 , n1418 ); 
nor ( n1420 , n1391 , n1419 ); 
nand ( n1421 , n1230 , n1242 ); 
nor ( n1422 , n1421 , n1258 ); 
buf ( n1423 , n1422 ); 
not ( n1424 , n1423 ); 
or ( n1425 , n1420 , n1424 ); 
nand ( n1426 , n1230 , n1251 ); 
not ( n1427 , n1426 ); 
not ( n1428 , n1422 ); 
not ( n1429 , n1428 ); 
or ( n1430 , n1427 , n1429 ); 
nand ( n1431 , n1156 , n1186 ); 
nand ( n1432 , n1430 , n1431 ); 
and ( n1433 , n1432 , n61 ); 
and ( n1434 , n1422 , n1192 ); 
not ( n1435 , n1434 ); 
not ( n1436 , n974 ); 
or ( n1437 , n1435 , n1436 ); 
not ( n1438 , n1426 ); 
nand ( n1439 , n1438 , n926 ); 
not ( n1440 , n35 ); 
and ( n1441 , n39 , n47 ); 
nand ( n1442 , n1441 , n51 ); 
nor ( n1443 , n1440 , n1442 ); 
and ( n1444 , n43 , n1443 ); 
and ( n1445 , n67 , n1444 ); 
or ( n1446 , n1445 , n63 ); 
nand ( n1447 , n1445 , n63 ); 
nand ( n1448 , n1446 , n1447 ); 
or ( n1449 , n1439 , n1448 ); 
nand ( n1450 , n1437 , n1449 ); 
nor ( n1451 , n1433 , n1450 ); 
nand ( n1452 , n1425 , n1451 ); 
not ( n1453 , n1187 ); 
nor ( n1454 , n1119 , n384 ); 
and ( n1455 , n1454 , n352 ); 
nand ( n1456 , n1455 , n401 ); 
nand ( n1457 , n1127 , n1406 ); 
nor ( n1458 , n1456 , n1457 ); 
not ( n1459 , n1458 ); 
nand ( n1460 , n1459 , n1406 ); 
and ( n1461 , n1460 , n503 ); 
not ( n1462 , n1460 ); 
and ( n1463 , n1462 , n504 ); 
nor ( n1464 , n1461 , n1463 ); 
or ( n1465 , n1464 , n1393 ); 
not ( n1466 , n1404 ); 
xnor ( n1467 , n1125 , n401 ); 
or ( n1468 , n1466 , n1467 ); 
nand ( n1469 , n1465 , n1468 ); 
not ( n1470 , n1469 ); 
or ( n1471 , n1453 , n1470 ); 
not ( n1472 , n465 ); 
not ( n1473 , n1472 ); 
not ( n1474 , n601 ); 
not ( n1475 , n686 ); 
nand ( n1476 , n678 , n1475 ); 
not ( n1477 , n1476 ); 
or ( n1478 , n1474 , n1477 ); 
not ( n1479 , n688 ); 
nand ( n1480 , n1478 , n1479 ); 
and ( n1481 , n1480 , n552 ); 
not ( n1482 , n386 ); 
nor ( n1483 , n1481 , n1482 ); 
nand ( n1484 , n1483 , n420 ); 
nand ( n1485 , n1484 , n424 ); 
not ( n1486 , n1485 ); 
or ( n1487 , n1473 , n1486 ); 
or ( n1488 , n1485 , n1472 ); 
nand ( n1489 , n1487 , n1488 ); 
nand ( n1490 , n1489 , n932 ); 
nand ( n1491 , n1471 , n1490 ); 
xor ( n1492 , n1355 , n1348 ); 
nand ( n1493 , n964 , n1492 ); 
not ( n1494 , n1174 ); 
buf ( n1495 , n458 ); 
xor ( n1496 , n1494 , n1495 ); 
and ( n1497 , n1496 , n1189 ); 
and ( n1498 , n1192 , n1495 ); 
nor ( n1499 , n1497 , n1498 ); 
nand ( n1500 , n1493 , n1499 ); 
or ( n1501 , n1491 , n1500 ); 
nand ( n1502 , n1501 , n1423 ); 
and ( n1503 , n1432 , n42 ); 
not ( n1504 , n1439 ); 
xor ( n1505 , n43 , n1443 ); 
and ( n1506 , n1504 , n1505 ); 
nor ( n1507 , n1503 , n1506 ); 
nand ( n1508 , n1502 , n1507 ); 
not ( n1509 , n1261 ); 
nor ( n1510 , n1096 , n764 ); 
not ( n1511 , n1510 ); 
nand ( n1512 , n1511 , n1098 ); 
and ( n1513 , n1088 , n1512 ); 
not ( n1514 , n1088 ); 
and ( n1515 , n1098 , n1134 ); 
nor ( n1516 , n1515 , n831 ); 
or ( n1517 , n1516 , n940 ); 
nand ( n1518 , n1517 , n1137 , n1138 ); 
and ( n1519 , n1514 , n1518 ); 
nor ( n1520 , n1513 , n1519 ); 
not ( n1521 , n1520 ); 
or ( n1522 , n1521 , n1155 ); 
or ( n1523 , n1191 , n818 ); 
nand ( n1524 , n1522 , n1523 ); 
and ( n1525 , n1047 , n838 ); 
not ( n1526 , n1047 ); 
and ( n1527 , n1526 , n839 ); 
nor ( n1528 , n1525 , n1527 ); 
not ( n1529 , n1528 ); 
not ( n1530 , n1078 ); 
or ( n1531 , n1529 , n1530 ); 
or ( n1532 , n1078 , n1528 ); 
nand ( n1533 , n1531 , n1532 ); 
nor ( n1534 , n1533 , n1198 ); 
nor ( n1535 , n1524 , n1534 ); 
nand ( n1536 , n1285 , n1159 ); 
and ( n1537 , n1536 , n819 ); 
not ( n1538 , n1536 ); 
and ( n1539 , n1538 , n818 ); 
nor ( n1540 , n1537 , n1539 ); 
nand ( n1541 , n1540 , n1189 ); 
and ( n1542 , n766 , n838 ); 
not ( n1543 , n766 ); 
and ( n1544 , n1543 , n839 ); 
nor ( n1545 , n1542 , n1544 ); 
not ( n1546 , n1307 ); 
not ( n1547 , n1546 ); 
not ( n1548 , n769 ); 
or ( n1549 , n1547 , n1548 ); 
buf ( n1550 , n874 ); 
nand ( n1551 , n1549 , n1550 ); 
xor ( n1552 , n1545 , n1551 ); 
nand ( n1553 , n1552 , n932 ); 
nand ( n1554 , n1535 , n1541 , n1553 ); 
not ( n1555 , n1554 ); 
or ( n1556 , n1509 , n1555 ); 
not ( n1557 , n1261 ); 
nand ( n1558 , n1557 , n84 ); 
nand ( n1559 , n1556 , n1558 ); 
not ( n1560 , n64 ); 
not ( n1561 , n1262 ); 
or ( n1562 , n1560 , n1561 ); 
or ( n1563 , n1191 , n1436 ); 
nand ( n1564 , n1563 , n1418 , n1412 ); 
nor ( n1565 , n1391 , n1564 ); 
or ( n1566 , n1565 , n1262 ); 
nand ( n1567 , n1562 , n1566 ); 
not ( n1568 , n68 ); 
not ( n1569 , n1262 ); 
or ( n1570 , n1568 , n1569 ); 
nand ( n1571 , n1361 , n1363 ); 
not ( n1572 , n1571 ); 
not ( n1573 , n1359 ); 
or ( n1574 , n1572 , n1573 ); 
or ( n1575 , n1359 , n1571 ); 
nand ( n1576 , n1574 , n1575 ); 
and ( n1577 , n1576 , n964 ); 
or ( n1578 , n1494 , n1495 ); 
buf ( n1579 , n543 ); 
nand ( n1580 , n1578 , n1579 ); 
and ( n1581 , n1580 , n1176 , n1189 ); 
nor ( n1582 , n1577 , n1581 ); 
not ( n1583 , n1191 ); 
not ( n1584 , n1579 ); 
not ( n1585 , n1584 ); 
and ( n1586 , n1583 , n1585 ); 
not ( n1587 , n1381 ); 
not ( n1588 , n1378 ); 
and ( n1589 , n1587 , n1588 ); 
and ( n1590 , n1380 , n691 ); 
and ( n1591 , n1377 , n548 ); 
nor ( n1592 , n1590 , n1591 ); 
nor ( n1593 , n1589 , n1592 ); 
and ( n1594 , n1593 , n932 ); 
nor ( n1595 , n1586 , n1594 ); 
nand ( n1596 , n1582 , n1595 ); 
or ( n1597 , n1466 , n1457 ); 
not ( n1598 , n504 ); 
not ( n1599 , n1458 ); 
or ( n1600 , n1598 , n1599 ); 
nand ( n1601 , n1600 , n1107 ); 
nand ( n1602 , n1601 , n1394 , n1398 ); 
nand ( n1603 , n1597 , n1602 ); 
nor ( n1604 , n1596 , n1603 ); 
or ( n1605 , n1604 , n1262 ); 
nand ( n1606 , n1570 , n1605 ); 
not ( n1607 , n44 ); 
not ( n1608 , n1261 ); 
not ( n1609 , n1608 ); 
or ( n1610 , n1607 , n1609 ); 
not ( n1611 , n1490 ); 
nor ( n1612 , n1611 , n1500 , n1469 ); 
not ( n1613 , n1261 ); 
or ( n1614 , n1612 , n1613 ); 
nand ( n1615 , n1610 , n1614 ); 
not ( n1616 , n1192 ); 
not ( n1617 , n1231 ); 
nand ( n1618 , n1617 , n1234 , n1241 ); 
and ( n1619 , n1257 , n1229 ); 
nand ( n1620 , n1618 , n1226 , n1254 , n1619 ); 
buf ( n1621 , n1620 ); 
not ( n1622 , n1621 ); 
not ( n1623 , n1622 ); 
or ( n1624 , n1616 , n1623 ); 
nand ( n1625 , n1624 , n1439 ); 
and ( n1626 , n1625 , n1495 ); 
buf ( n1627 , n1188 ); 
not ( n1628 , n1627 ); 
not ( n1629 , n1620 ); 
nand ( n1630 , n1628 , n1629 ); 
not ( n1631 , n1630 ); 
and ( n1632 , n1631 , n1496 ); 
and ( n1633 , n1228 , n43 ); 
nor ( n1634 , n1626 , n1632 , n1633 ); 
nand ( n1635 , n1629 , n1192 ); 
and ( n1636 , n1439 , n1635 ); 
not ( n1637 , n928 ); 
nand ( n1638 , n923 , n1187 ); 
not ( n1639 , n1638 ); 
or ( n1640 , n1637 , n1639 ); 
nand ( n1641 , n1640 , n1629 ); 
and ( n1642 , n1641 , n1630 , n158 ); 
nand ( n1643 , n1636 , n1642 ); 
not ( n1644 , n1643 ); 
nand ( n1645 , n1505 , n1644 ); 
not ( n1646 , n1493 ); 
or ( n1647 , n1491 , n1646 ); 
not ( n1648 , n1622 ); 
buf ( n1649 , n1648 ); 
buf ( n1650 , n1649 ); 
not ( n1651 , n1650 ); 
nand ( n1652 , n1647 , n1651 ); 
nand ( n1653 , n1634 , n1645 , n1652 ); 
not ( n1654 , n1286 ); 
or ( n1655 , n1285 , n1158 ); 
nand ( n1656 , n1655 , n1189 ); 
not ( n1657 , n1656 ); 
and ( n1658 , n1654 , n1657 ); 
not ( n1659 , n1273 ); 
nand ( n1660 , n1072 , n968 ); 
not ( n1661 , n1660 ); 
or ( n1662 , n1659 , n1661 ); 
or ( n1663 , n1273 , n1660 ); 
nand ( n1664 , n1662 , n1663 ); 
and ( n1665 , n964 , n1664 ); 
nor ( n1666 , n1658 , n1665 ); 
not ( n1667 , n1311 ); 
nand ( n1668 , n1667 , n1300 ); 
and ( n1669 , n1300 , n1310 ); 
nor ( n1670 , n1669 , n1303 ); 
and ( n1671 , n1307 , n1670 ); 
nor ( n1672 , n1671 , n933 ); 
and ( n1673 , n1668 , n1672 ); 
nor ( n1674 , n1158 , n1191 ); 
nor ( n1675 , n1673 , n1674 ); 
nand ( n1676 , n1666 , n1675 ); 
not ( n1677 , n1315 ); 
and ( n1678 , n1512 , n1131 ); 
nor ( n1679 , n1678 , n1393 ); 
not ( n1680 , n1679 ); 
or ( n1681 , n1677 , n1680 ); 
and ( n1682 , n797 , n1395 ); 
or ( n1683 , n1682 , n702 ); 
nand ( n1684 , n1683 , n1324 ); 
or ( n1685 , n1466 , n1684 ); 
nand ( n1686 , n1681 , n1685 ); 
nor ( n1687 , n1676 , n1686 ); 
or ( n1688 , n1687 , n1262 ); 
not ( n1689 , n72 ); 
or ( n1690 , n1689 , n1261 ); 
nand ( n1691 , n1688 , n1690 ); 
or ( n1692 , n1687 , n1339 ); 
not ( n1693 , n70 ); 
or ( n1694 , n1693 , n1338 ); 
nand ( n1695 , n1692 , n1694 ); 
not ( n1696 , n62 ); 
not ( n1697 , n1339 ); 
or ( n1698 , n1696 , n1697 ); 
or ( n1699 , n1565 , n1339 ); 
nand ( n1700 , n1698 , n1699 ); 
not ( n1701 , n66 ); 
not ( n1702 , n1339 ); 
or ( n1703 , n1701 , n1702 ); 
or ( n1704 , n1604 , n1339 ); 
nand ( n1705 , n1703 , n1704 ); 
not ( n1706 , n41 ); 
not ( n1707 , n1339 ); 
or ( n1708 , n1706 , n1707 ); 
or ( n1709 , n1612 , n1339 ); 
nand ( n1710 , n1708 , n1709 ); 
not ( n1711 , n54 ); 
not ( n1712 , n1339 ); 
or ( n1713 , n1711 , n1712 ); 
not ( n1714 , n804 ); 
and ( n1715 , n550 , n691 ); 
not ( n1716 , n1715 ); 
or ( n1717 , n1714 , n1716 ); 
nand ( n1718 , n1717 , n856 ); 
and ( n1719 , n798 , n777 ); 
not ( n1720 , n798 ); 
and ( n1721 , n1720 , n776 ); 
nor ( n1722 , n1719 , n1721 ); 
xor ( n1723 , n1718 , n1722 ); 
nand ( n1724 , n1723 , n932 ); 
not ( n1725 , n976 ); 
not ( n1726 , n1062 ); 
not ( n1727 , n1039 ); 
or ( n1728 , n1726 , n1727 ); 
not ( n1729 , n1041 ); 
nand ( n1730 , n1728 , n1729 ); 
not ( n1731 , n1730 ); 
or ( n1732 , n1725 , n1731 ); 
not ( n1733 , n975 ); 
not ( n1734 , n1042 ); 
or ( n1735 , n1733 , n1734 ); 
nand ( n1736 , n1735 , n855 ); 
nand ( n1737 , n1732 , n1736 ); 
not ( n1738 , n1737 ); 
nand ( n1739 , n1069 , n982 ); 
not ( n1740 , n1739 ); 
nor ( n1741 , n1198 , n1740 ); 
nand ( n1742 , n1738 , n1741 ); 
nor ( n1743 , n1198 , n1739 ); 
and ( n1744 , n1737 , n1743 ); 
not ( n1745 , n774 ); 
not ( n1746 , n1192 ); 
or ( n1747 , n1745 , n1746 ); 
not ( n1748 , n1285 ); 
not ( n1749 , n1284 ); 
not ( n1750 , n1161 ); 
and ( n1751 , n1749 , n1750 ); 
nor ( n1752 , n1751 , n1416 ); 
nand ( n1753 , n1748 , n1752 ); 
nand ( n1754 , n1747 , n1753 ); 
nor ( n1755 , n1744 , n1754 ); 
nand ( n1756 , n1724 , n1742 , n1755 ); 
not ( n1757 , n969 ); 
not ( n1758 , n1130 ); 
nand ( n1759 , n1324 , n1758 ); 
not ( n1760 , n1759 ); 
or ( n1761 , n1757 , n1760 ); 
or ( n1762 , n1759 , n969 ); 
nand ( n1763 , n1761 , n1762 ); 
and ( n1764 , n1763 , n1394 ); 
and ( n1765 , n1404 , n1396 ); 
nor ( n1766 , n1764 , n1765 ); 
not ( n1767 , n1766 ); 
nor ( n1768 , n1756 , n1767 ); 
or ( n1769 , n1768 , n1339 ); 
nand ( n1770 , n1713 , n1769 ); 
or ( n1771 , n1420 , n1650 ); 
not ( n1772 , n1448 ); 
and ( n1773 , n1644 , n1772 ); 
not ( n1774 , n63 ); 
not ( n1775 , n1228 ); 
or ( n1776 , n1774 , n1775 ); 
buf ( n1777 , n1636 ); 
or ( n1778 , n1777 , n1436 ); 
nand ( n1779 , n1776 , n1778 ); 
nor ( n1780 , n1773 , n1779 ); 
nand ( n1781 , n1771 , n1780 ); 
not ( n1782 , n1338 ); 
not ( n1783 , n1554 ); 
or ( n1784 , n1782 , n1783 ); 
nand ( n1785 , n1339 , n82 ); 
nand ( n1786 , n1784 , n1785 ); 
not ( n1787 , n1596 ); 
or ( n1788 , n1787 , n1424 ); 
and ( n1789 , n1432 , n65 ); 
and ( n1790 , n1422 , n1187 ); 
and ( n1791 , n1790 , n1603 ); 
xor ( n1792 , n67 , n1444 ); 
and ( n1793 , n1504 , n1792 ); 
nor ( n1794 , n1789 , n1791 , n1793 ); 
nand ( n1795 , n1788 , n1794 ); 
not ( n1796 , n1676 ); 
or ( n1797 , n1796 , n1424 ); 
and ( n1798 , n1432 , n69 ); 
not ( n1799 , n1447 ); 
and ( n1800 , n57 , n1799 ); 
nand ( n1801 , n1800 , n55 ); 
not ( n1802 , n1801 ); 
xor ( n1803 , n71 , n1802 ); 
and ( n1804 , n1504 , n1803 ); 
and ( n1805 , n1790 , n1686 ); 
nor ( n1806 , n1798 , n1804 , n1805 ); 
nand ( n1807 , n1797 , n1806 ); 
not ( n1808 , n1715 ); 
nand ( n1809 , n1365 , n851 ); 
nand ( n1810 , n1808 , n1809 ); 
not ( n1811 , n855 ); 
and ( n1812 , n803 , n1811 ); 
not ( n1813 , n803 ); 
and ( n1814 , n1813 , n855 ); 
nor ( n1815 , n1812 , n1814 ); 
nor ( n1816 , n1810 , n1815 ); 
not ( n1817 , n1816 ); 
nand ( n1818 , n1810 , n1815 ); 
nand ( n1819 , n1817 , n1818 , n932 ); 
and ( n1820 , n1811 , n975 ); 
not ( n1821 , n1811 ); 
and ( n1822 , n1821 , n976 ); 
nor ( n1823 , n1820 , n1822 ); 
not ( n1824 , n1730 ); 
xor ( n1825 , n1823 , n1824 ); 
and ( n1826 , n1825 , n964 ); 
or ( n1827 , n1178 , n1160 ); 
nand ( n1828 , n1827 , n1189 ); 
nor ( n1829 , n1284 , n1828 ); 
nor ( n1830 , n1826 , n1829 ); 
not ( n1831 , n1398 ); 
nand ( n1832 , n1831 , n797 ); 
and ( n1833 , n1832 , n1684 ); 
nor ( n1834 , n1833 , n1393 ); 
and ( n1835 , n1834 , n1758 ); 
not ( n1836 , n1107 ); 
and ( n1837 , n1404 , n1836 ); 
nor ( n1838 , n1835 , n1837 ); 
nand ( n1839 , n1819 , n1830 , n1838 ); 
nand ( n1840 , n1819 , n1830 , n1186 ); 
nand ( n1841 , n1839 , n1840 ); 
or ( n1842 , n1841 , n1424 ); 
and ( n1843 , n1432 , n58 ); 
xor ( n1844 , n57 , n1799 ); 
not ( n1845 , n1844 ); 
not ( n1846 , n1504 ); 
or ( n1847 , n1845 , n1846 ); 
or ( n1848 , n1435 , n1160 ); 
nand ( n1849 , n1847 , n1848 ); 
nor ( n1850 , n1843 , n1849 ); 
nand ( n1851 , n1842 , n1850 ); 
not ( n1852 , n60 ); 
not ( n1853 , n1262 ); 
or ( n1854 , n1852 , n1853 ); 
nor ( n1855 , n1191 , n1160 ); 
nor ( n1856 , n1839 , n1855 ); 
or ( n1857 , n1856 , n1262 ); 
nand ( n1858 , n1854 , n1857 ); 
not ( n1859 , n36 ); 
not ( n1860 , n1262 ); 
or ( n1861 , n1859 , n1860 ); 
not ( n1862 , n1168 ); 
and ( n1863 , n1192 , n1862 ); 
not ( n1864 , n1484 ); 
or ( n1865 , n1483 , n420 ); 
nand ( n1866 , n1865 , n931 ); 
nor ( n1867 , n1864 , n1866 ); 
not ( n1868 , n1867 ); 
and ( n1869 , n1017 , n1025 ); 
not ( n1870 , n1353 ); 
and ( n1871 , n1869 , n1870 ); 
nor ( n1872 , n1871 , n1197 ); 
buf ( n1873 , n1354 ); 
and ( n1874 , n1872 , n1873 ); 
nor ( n1875 , n1170 , n675 ); 
nand ( n1876 , n1875 , n1172 ); 
nor ( n1877 , n1876 , n1165 ); 
not ( n1878 , n1877 ); 
nand ( n1879 , n1878 , n1862 ); 
and ( n1880 , n1494 , n1879 , n1189 ); 
nor ( n1881 , n1874 , n1880 ); 
and ( n1882 , n1456 , n1457 ); 
nor ( n1883 , n1882 , n1458 ); 
and ( n1884 , n1394 , n1883 ); 
not ( n1885 , n1124 ); 
or ( n1886 , n1885 , n352 ); 
not ( n1887 , n1125 ); 
nand ( n1888 , n1886 , n1887 ); 
not ( n1889 , n1888 ); 
and ( n1890 , n1404 , n1889 ); 
nor ( n1891 , n1884 , n1890 ); 
and ( n1892 , n1868 , n1881 , n1891 ); 
not ( n1893 , n1892 ); 
nor ( n1894 , n1863 , n1893 ); 
or ( n1895 , n1894 , n1613 ); 
nand ( n1896 , n1861 , n1895 ); 
not ( n1897 , n59 ); 
not ( n1898 , n1339 ); 
or ( n1899 , n1897 , n1898 ); 
or ( n1900 , n1856 , n1339 ); 
nand ( n1901 , n1899 , n1900 ); 
not ( n1902 , n1582 ); 
and ( n1903 , n1603 , n1187 ); 
nor ( n1904 , n1902 , n1903 ); 
or ( n1905 , n1904 , n1650 ); 
and ( n1906 , n1644 , n1792 ); 
not ( n1907 , n1593 ); 
and ( n1908 , n1622 , n931 ); 
not ( n1909 , n1908 ); 
or ( n1910 , n1907 , n1909 ); 
or ( n1911 , n1777 , n1584 ); 
not ( n1912 , n67 ); 
or ( n1913 , n1912 , n158 ); 
nand ( n1914 , n1910 , n1911 , n1913 ); 
nor ( n1915 , n1906 , n1914 ); 
nand ( n1916 , n1905 , n1915 ); 
or ( n1917 , n1841 , n1650 ); 
and ( n1918 , n1644 , n1844 ); 
or ( n1919 , n1777 , n1160 ); 
not ( n1920 , n57 ); 
or ( n1921 , n1920 , n158 ); 
nand ( n1922 , n1919 , n1921 ); 
nor ( n1923 , n1918 , n1922 ); 
nand ( n1924 , n1917 , n1923 ); 
or ( n1925 , n1650 , n1293 ); 
not ( n1926 , n1909 ); 
nand ( n1927 , n1926 , n1312 ); 
not ( n1928 , n1777 ); 
and ( n1929 , n71 , n1802 ); 
or ( n1930 , n1929 , n75 ); 
nand ( n1931 , n1929 , n75 ); 
nand ( n1932 , n1930 , n1931 ); 
not ( n1933 , n1932 ); 
nand ( n1934 , n1933 , n1642 ); 
not ( n1935 , n1934 ); 
or ( n1936 , n1928 , n1935 ); 
or ( n1937 , n1777 , n1046 ); 
nand ( n1938 , n1936 , n1937 ); 
nor ( n1939 , n1648 , n1638 ); 
and ( n1940 , n1328 , n1939 ); 
and ( n1941 , n1228 , n75 ); 
nor ( n1942 , n1940 , n1941 ); 
and ( n1943 , n1927 , n1938 , n1942 ); 
nand ( n1944 , n1925 , n1943 ); 
not ( n1945 , n1442 ); 
not ( n1946 , n35 ); 
and ( n1947 , n1945 , n1946 ); 
and ( n1948 , n1442 , n35 ); 
nor ( n1949 , n1947 , n1948 ); 
or ( n1950 , n1643 , n1949 ); 
not ( n1951 , n1881 ); 
nor ( n1952 , n1951 , n1187 , n1867 ); 
nor ( n1953 , n1952 , n1892 ); 
nand ( n1954 , n1953 , n1651 ); 
and ( n1955 , n1625 , n1862 ); 
and ( n1956 , n1228 , n35 ); 
nor ( n1957 , n1955 , n1956 ); 
nand ( n1958 , n1950 , n1954 , n1957 ); 
not ( n1959 , n34 ); 
not ( n1960 , n1339 ); 
or ( n1961 , n1959 , n1960 ); 
or ( n1962 , n1894 , n1339 ); 
nand ( n1963 , n1961 , n1962 ); 
not ( n1964 , n1534 ); 
not ( n1965 , n1964 ); 
not ( n1966 , n1541 ); 
or ( n1967 , n1965 , n1966 ); 
nand ( n1968 , n1967 , n1651 ); 
not ( n1969 , n1931 ); 
or ( n1970 , n1969 , n83 ); 
nand ( n1971 , n1969 , n83 ); 
nand ( n1972 , n1970 , n1644 , n1971 ); 
and ( n1973 , n1552 , n1908 ); 
or ( n1974 , n1777 , n818 ); 
and ( n1975 , n1520 , n1939 ); 
and ( n1976 , n1228 , n83 ); 
nor ( n1977 , n1975 , n1976 ); 
nand ( n1978 , n1974 , n1977 ); 
nor ( n1979 , n1973 , n1978 ); 
nand ( n1980 , n1968 , n1972 , n1979 ); 
not ( n1981 , n1423 ); 
not ( n1982 , n1953 ); 
or ( n1983 , n1981 , n1982 ); 
and ( n1984 , n1432 , n33 ); 
or ( n1985 , n1435 , n1168 ); 
or ( n1986 , n1439 , n1949 ); 
nand ( n1987 , n1985 , n1986 ); 
nor ( n1988 , n1984 , n1987 ); 
nand ( n1989 , n1983 , n1988 ); 
not ( n1990 , n1423 ); 
not ( n1991 , n1756 ); 
or ( n1992 , n1990 , n1991 ); 
and ( n1993 , n1432 , n53 ); 
and ( n1994 , n1790 , n1767 ); 
or ( n1995 , n1800 , n55 ); 
nand ( n1996 , n1995 , n1801 ); 
nor ( n1997 , n1439 , n1996 ); 
nor ( n1998 , n1993 , n1994 , n1997 ); 
nand ( n1999 , n1992 , n1998 ); 
and ( n2000 , n1737 , n1739 ); 
not ( n2001 , n1737 ); 
and ( n2002 , n2001 , n1740 ); 
nor ( n2003 , n2000 , n2002 ); 
and ( n2004 , n2003 , n964 ); 
not ( n2005 , n1753 ); 
nor ( n2006 , n2004 , n2005 ); 
or ( n2007 , n2006 , n1650 ); 
not ( n2008 , n1643 ); 
not ( n2009 , n1996 ); 
and ( n2010 , n2008 , n2009 ); 
not ( n2011 , n1723 ); 
or ( n2012 , n2011 , n1909 ); 
and ( n2013 , n1625 , n774 ); 
not ( n2014 , n1621 ); 
nand ( n2015 , n2014 , n1187 ); 
or ( n2016 , n2015 , n1766 ); 
or ( n2017 , n697 , n158 ); 
nand ( n2018 , n2016 , n2017 ); 
nor ( n2019 , n2013 , n2018 ); 
nand ( n2020 , n2012 , n2019 ); 
nor ( n2021 , n2010 , n2020 ); 
nand ( n2022 , n2007 , n2021 ); 
not ( n2023 , n879 ); 
and ( n2024 , n956 , n2023 ); 
not ( n2025 , n956 ); 
and ( n2026 , n2025 , n879 ); 
nor ( n2027 , n2024 , n2026 ); 
nor ( n2028 , n2027 , n1909 ); 
not ( n2029 , n1971 ); 
not ( n2030 , n77 ); 
and ( n2031 , n2029 , n2030 ); 
and ( n2032 , n1971 , n77 ); 
nor ( n2033 , n2031 , n2032 ); 
nor ( n2034 , n2033 , n1643 ); 
and ( n2035 , n1625 , n950 ); 
and ( n2036 , n1228 , n77 ); 
nor ( n2037 , n2035 , n2036 ); 
and ( n2038 , n1153 , n1939 ); 
and ( n2039 , n1183 , n1631 ); 
nor ( n2040 , n2038 , n2039 ); 
nand ( n2041 , n2037 , n2040 ); 
nor ( n2042 , n2028 , n2034 , n2041 ); 
not ( n2043 , n1666 ); 
nand ( n2044 , n2043 , n1651 ); 
and ( n2045 , n1644 , n1803 ); 
not ( n2046 , n1668 ); 
not ( n2047 , n1671 ); 
nand ( n2048 , n2047 , n1908 ); 
or ( n2049 , n2046 , n2048 ); 
not ( n2050 , n71 ); 
not ( n2051 , n1228 ); 
or ( n2052 , n2050 , n2051 ); 
or ( n2053 , n1777 , n1158 ); 
nand ( n2054 , n2052 , n2053 ); 
not ( n2055 , n1686 ); 
nor ( n2056 , n2055 , n2015 ); 
nor ( n2057 , n2054 , n2056 ); 
nand ( n2058 , n2049 , n2057 ); 
nor ( n2059 , n2045 , n2058 ); 
nand ( n2060 , n2044 , n2059 ); 
or ( n2061 , n1196 , n965 ); 
nand ( n2062 , n2061 , n1200 ); 
or ( n2063 , n1643 , n39 ); 
not ( n2064 , n1172 ); 
and ( n2065 , n1625 , n2064 ); 
not ( n2066 , n1638 ); 
buf ( n2067 , n1475 ); 
not ( n2068 , n2067 ); 
nand ( n2069 , n2068 , n679 ); 
nand ( n2070 , n2069 , n929 , n1476 ); 
not ( n2071 , n1005 ); 
buf ( n2072 , n1008 ); 
or ( n2073 , n1875 , n1172 ); 
not ( n2074 , n1188 ); 
nand ( n2075 , n2073 , n2074 , n1876 ); 
and ( n2076 , n2070 , t_0 , n2075 ); 
not ( n2077 , n2076 ); 
or ( n2078 , n2066 , n2077 ); 
not ( n2079 , n1009 ); 
and ( n2080 , n1119 , n384 , n2079 ); 
not ( n2081 , n1885 ); 
nand ( n2082 , n2081 , n1321 ); 
nor ( n2083 , n2080 , n2082 ); 
not ( n2084 , n1454 ); 
and ( n2085 , n2083 , n2084 ); 
and ( n2086 , n1088 , n611 ); 
nor ( n2087 , n2085 , n2086 ); 
nand ( n2088 , n2076 , n2087 ); 
nand ( n2089 , n2078 , n2088 ); 
or ( n2090 , n1649 , n2089 ); 
not ( n2091 , n39 ); 
or ( n2092 , n2091 , n158 ); 
nand ( n2093 , n2090 , n2092 ); 
nor ( n2094 , n2065 , n2093 ); 
nand ( n2095 , n2063 , n2094 ); 
or ( n2096 , n1441 , n51 ); 
nand ( n2097 , n2096 , n1442 ); 
or ( n2098 , n1643 , n2097 ); 
buf ( n2099 , n357 ); 
xor ( n2100 , n385 , n2099 ); 
xnor ( n2101 , n2100 , n690 ); 
nand ( n2102 , n2101 , n931 ); 
buf ( n2103 , n1017 ); 
buf ( n2104 , n1010 ); 
not ( n2105 , n2104 ); 
not ( n2106 , n556 ); 
not ( n2107 , n2106 ); 
and ( n2108 , n2105 , n2107 ); 
and ( n2109 , n2106 , n2104 ); 
nor ( n2110 , n2108 , n2109 ); 
or ( n2111 , n2110 , n2072 ); 
nand ( n2112 , n2111 , n1014 , n1011 ); 
and ( n2113 , n2103 , n2112 , n963 ); 
not ( n2114 , n1876 ); 
buf ( n2115 , n1164 ); 
and ( n2116 , n2114 , n2115 ); 
buf ( n2117 , n388 ); 
nor ( n2118 , n2116 , n2117 ); 
nor ( n2119 , n1188 , n2118 , n1877 ); 
nor ( n2120 , n2113 , n2119 ); 
nand ( n2121 , n2102 , n1186 , n2120 ); 
not ( n2122 , n1455 ); 
and ( n2123 , n2122 , n1467 ); 
not ( n2124 , n2122 ); 
and ( n2125 , n2124 , n401 ); 
nor ( n2126 , n2123 , n2125 ); 
and ( n2127 , n1394 , n2126 ); 
and ( n2128 , n384 , n2079 ); 
not ( n2129 , n384 ); 
and ( n2130 , n2129 , n1009 ); 
nor ( n2131 , n2128 , n2130 ); 
and ( n2132 , n1404 , n2131 ); 
nor ( n2133 , n2127 , n2132 ); 
nand ( n2134 , n2120 , n2102 , n2133 ); 
not ( n2135 , n1648 ); 
nand ( n2136 , n2121 , n2134 , n2135 ); 
not ( n2137 , n2117 ); 
nand ( n2138 , n1625 , n2137 ); 
nand ( n2139 , n1228 , n51 ); 
and ( n2140 , n2136 , n2138 , n2139 ); 
nand ( n2141 , n2098 , n2140 ); 
not ( n2142 , n2089 ); 
nand ( n2143 , n2142 , n1423 ); 
nand ( n2144 , n1434 , n2064 ); 
nand ( n2145 , n1432 , n37 ); 
nand ( n2146 , n2091 , n1504 ); 
nand ( n2147 , n2143 , n2144 , n2145 , n2146 ); 
nand ( n2148 , n2121 , n2134 , n1423 ); 
nand ( n2149 , n1434 , n2137 ); 
nand ( n2150 , n1432 , n49 ); 
not ( n2151 , n2097 ); 
nand ( n2152 , n2151 , n1504 ); 
nand ( n2153 , n2148 , n2149 , n2150 , n2152 ); 
not ( n2154 , n154 ); 
nand ( n2155 , n1643 , n158 ); 
not ( n2156 , n2155 ); 
or ( n2157 , n2154 , n2156 ); 
and ( n2158 , n1625 , n675 ); 
not ( n2159 , n1908 ); 
not ( n2160 , n672 ); 
nor ( n2161 , n2160 , n639 ); 
not ( n2162 , n2161 ); 
not ( n2163 , n618 ); 
nand ( n2164 , n2163 , n677 ); 
not ( n2165 , n2164 ); 
or ( n2166 , n2162 , n2165 ); 
or ( n2167 , n2161 , n2164 ); 
nand ( n2168 , n2166 , n2167 ); 
not ( n2169 , n2168 ); 
or ( n2170 , n2159 , n2169 ); 
not ( n2171 , n1649 ); 
not ( n2172 , n987 ); 
nand ( n2173 , n2172 , n2071 , n997 ); 
not ( n2174 , n2173 ); 
not ( n2175 , n2164 ); 
or ( n2176 , n2174 , n2175 ); 
or ( n2177 , n2173 , n2164 ); 
nand ( n2178 , n2176 , n2177 ); 
and ( n2179 , n963 , n2178 ); 
and ( n2180 , n1170 , n675 ); 
nor ( n2181 , n2180 , n1875 , n1188 ); 
nor ( n2182 , n2179 , n2181 ); 
not ( n2183 , n2182 ); 
and ( n2184 , n2171 , n2183 ); 
not ( n2185 , n2015 ); 
not ( n2186 , n636 ); 
not ( n2187 , n1404 ); 
or ( n2188 , n2186 , n2187 ); 
not ( n2189 , n1117 ); 
or ( n2190 , n2189 , n610 ); 
nand ( n2191 , n2190 , n598 ); 
nand ( n2192 , n1394 , n2191 , n1119 ); 
nand ( n2193 , n2188 , n2192 ); 
and ( n2194 , n2185 , n2193 ); 
nor ( n2195 , n2184 , n2194 ); 
nand ( n2196 , n2170 , n2195 ); 
nor ( n2197 , n2158 , n2196 ); 
nand ( n2198 , n2157 , n2197 ); 
not ( n2199 , n146 ); 
not ( n2200 , n2155 ); 
or ( n2201 , n2199 , n2200 ); 
nand ( n2202 , n1777 , n1630 ); 
buf ( n2203 , n658 ); 
not ( n2204 , n2203 ); 
and ( n2205 , n2202 , n2204 ); 
and ( n2206 , n2203 , n670 ); 
nor ( n2207 , n2206 , n671 ); 
nor ( n2208 , n928 , n2207 ); 
not ( n2209 , n2208 ); 
not ( n2210 , n2135 ); 
or ( n2211 , n2209 , n2210 ); 
or ( n2212 , n636 , n1116 ); 
nand ( n2213 , n2212 , n1394 , n2189 ); 
or ( n2214 , n2015 , n2213 ); 
nand ( n2215 , n2211 , n2214 ); 
nor ( n2216 , n2205 , n2215 ); 
nand ( n2217 , n2201 , n2216 ); 
and ( n2218 , n377 , n39 ); 
and ( n2219 , n2091 , n47 ); 
nor ( n2220 , n2218 , n2219 ); 
or ( n2221 , n1643 , n2220 ); 
not ( n2222 , n2115 ); 
and ( n2223 , n1625 , n2222 ); 
not ( n2224 , n1466 ); 
not ( n2225 , n598 ); 
and ( n2226 , n2224 , n2225 ); 
and ( n2227 , n2084 , n1888 ); 
nor ( n2228 , n2227 , n1455 , n1393 ); 
nor ( n2229 , n2226 , n2228 ); 
or ( n2230 , n2015 , n2229 ); 
not ( n2231 , n1476 ); 
not ( n2232 , n601 ); 
nor ( n2233 , n2232 , n688 ); 
not ( n2234 , n2233 ); 
or ( n2235 , n2231 , n2234 ); 
or ( n2236 , n1476 , n2233 ); 
nand ( n2237 , n2235 , n2236 ); 
not ( n2238 , n2237 ); 
not ( n2239 , n931 ); 
or ( n2240 , n2238 , n2239 ); 
xor ( n2241 , n2072 , n2110 ); 
and ( n2242 , n2241 , n963 ); 
not ( n2243 , n1188 ); 
not ( n2244 , n2222 ); 
not ( n2245 , n2114 ); 
or ( n2246 , n2244 , n2245 ); 
or ( n2247 , n2114 , n2222 ); 
nand ( n2248 , n2246 , n2247 ); 
and ( n2249 , n2243 , n2248 ); 
nor ( n2250 , n2242 , n2249 ); 
nand ( n2251 , n2240 , n2250 ); 
and ( n2252 , n2251 , n2135 ); 
and ( n2253 , n1228 , n47 ); 
nor ( n2254 , n2252 , n2253 ); 
nand ( n2255 , n2230 , n2254 ); 
nor ( n2256 , n2223 , n2255 ); 
nand ( n2257 , n2221 , n2256 ); 
not ( n2258 , n40 ); 
not ( n2259 , n1557 ); 
or ( n2260 , n2258 , n2259 ); 
nand ( n2261 , n2076 , n1155 ); 
and ( n2262 , n2088 , n2261 ); 
and ( n2263 , n1192 , n2064 ); 
nor ( n2264 , n2262 , n2263 ); 
or ( n2265 , n2264 , n1262 ); 
nand ( n2266 , n2260 , n2265 ); 
not ( n2267 , n150 ); 
not ( n2268 , n2155 ); 
or ( n2269 , n2267 , n2268 ); 
not ( n2270 , n648 ); 
and ( n2271 , n1625 , n2270 ); 
xnor ( n2272 , n2189 , n611 ); 
and ( n2273 , n1394 , n2272 ); 
and ( n2274 , n1404 , n670 ); 
nor ( n2275 , n2273 , n2274 ); 
or ( n2276 , n2015 , n2275 ); 
not ( n2277 , n1648 ); 
not ( n2278 , n1197 ); 
buf ( n2279 , n652 ); 
not ( n2280 , n2279 ); 
not ( n2281 , n986 ); 
and ( n2282 , n2280 , n2281 ); 
and ( n2283 , n2279 , n986 ); 
nor ( n2284 , n2282 , n2283 ); 
not ( n2285 , n2284 ); 
and ( n2286 , n2278 , n2285 ); 
or ( n2287 , n2279 , n671 ); 
nand ( n2288 , n2287 , n672 ); 
not ( n2289 , n2288 ); 
nor ( n2290 , n2289 , n930 ); 
nor ( n2291 , n2286 , n2290 ); 
not ( n2292 , n2291 ); 
and ( n2293 , n2277 , n2292 ); 
not ( n2294 , n2270 ); 
or ( n2295 , n2294 , n2203 ); 
nand ( n2296 , n2295 , n1170 ); 
nor ( n2297 , n1630 , n2296 ); 
nor ( n2298 , n2293 , n2297 ); 
nand ( n2299 , n2276 , n2298 ); 
nor ( n2300 , n2271 , n2299 ); 
nand ( n2301 , n2269 , n2300 ); 
not ( n2302 , n1339 ); 
not ( n2303 , n38 ); 
or ( n2304 , n2302 , n2303 ); 
or ( n2305 , n2264 , n1339 ); 
nand ( n2306 , n2304 , n2305 ); 
not ( n2307 , n52 ); 
not ( n2308 , n1608 ); 
or ( n2309 , n2307 , n2308 ); 
and ( n2310 , n1192 , n2137 ); 
nor ( n2311 , n2310 , n2134 ); 
or ( n2312 , n2311 , n1262 ); 
nand ( n2313 , n2309 , n2312 ); 
not ( n2314 , n1191 ); 
not ( n2315 , n2115 ); 
and ( n2316 , n2314 , n2315 ); 
nor ( n2317 , n2316 , n2251 ); 
not ( n2318 , n2317 ); 
nand ( n2319 , n2318 , n1423 ); 
not ( n2320 , n2229 ); 
and ( n2321 , n2320 , n1790 ); 
not ( n2322 , n2220 ); 
and ( n2323 , n1504 , n2322 ); 
nor ( n2324 , n2321 , n2323 ); 
nand ( n2325 , n1432 , n48 ); 
nand ( n2326 , n2319 , n2324 , n2325 ); 
not ( n2327 , n1339 ); 
not ( n2328 , n50 ); 
or ( n2329 , n2327 , n2328 ); 
or ( n2330 , n2311 , n1339 ); 
nand ( n2331 , n2329 , n2330 ); 
not ( n2332 , n155 ); 
not ( n2333 , n1432 ); 
or ( n2334 , n2332 , n2333 ); 
and ( n2335 , n154 , n1504 ); 
not ( n2336 , n1428 ); 
and ( n2337 , n931 , n2168 ); 
and ( n2338 , n1192 , n675 ); 
nor ( n2339 , n2337 , n2338 ); 
nand ( n2340 , n2182 , n2339 ); 
and ( n2341 , n2336 , n2340 ); 
not ( n2342 , n2193 ); 
not ( n2343 , n1790 ); 
nor ( n2344 , n2342 , n2343 ); 
nor ( n2345 , n2335 , n2341 , n2344 ); 
nand ( n2346 , n2334 , n2345 ); 
not ( n2347 , n1339 ); 
not ( n2348 , n46 ); 
or ( n2349 , n2347 , n2348 ); 
and ( n2350 , n2317 , n2229 ); 
or ( n2351 , n2350 , n1339 ); 
nand ( n2352 , n2349 , n2351 ); 
not ( n2353 , n147 ); 
not ( n2354 , n1432 ); 
or ( n2355 , n2353 , n2354 ); 
nor ( n2356 , n2343 , n2213 ); 
not ( n2357 , n146 ); 
not ( n2358 , n1504 ); 
or ( n2359 , n2357 , n2358 ); 
nand ( n2360 , n1188 , n1191 ); 
and ( n2361 , n2360 , n2204 ); 
nor ( n2362 , n2361 , n2208 ); 
not ( n2363 , n2362 ); 
nand ( n2364 , n2363 , n2336 ); 
nand ( n2365 , n2359 , n2364 ); 
nor ( n2366 , n2356 , n2365 ); 
nand ( n2367 , n2355 , n2366 ); 
not ( n2368 , n45 ); 
not ( n2369 , n1608 ); 
or ( n2370 , n2368 , n2369 ); 
or ( n2371 , n2350 , n1613 ); 
nand ( n2372 , n2370 , n2371 ); 
not ( n2373 , n153 ); 
not ( n2374 , n1432 ); 
or ( n2375 , n2373 , n2374 ); 
and ( n2376 , n150 , n1504 ); 
or ( n2377 , n1627 , n2296 ); 
or ( n2378 , n1191 , n2294 ); 
nand ( n2379 , n2377 , n2378 ); 
not ( n2380 , n2379 ); 
nand ( n2381 , n2380 , n2291 ); 
and ( n2382 , n2336 , n2381 ); 
nor ( n2383 , n2343 , n2275 ); 
nor ( n2384 , n2376 , n2382 , n2383 ); 
nand ( n2385 , n2375 , n2384 ); 
nor ( n2386 , n2340 , n2193 ); 
or ( n2387 , n2386 , n1262 ); 
nand ( n2388 , n1557 , n156 ); 
nand ( n2389 , n2387 , n2388 ); 
or ( n2390 , n2386 , n1339 ); 
nand ( n2391 , n1339 , n157 ); 
nand ( n2392 , n2390 , n2391 ); 
not ( n2393 , n2275 ); 
nor ( n2394 , n2393 , n2381 ); 
or ( n2395 , n1339 , n2394 ); 
nand ( n2396 , n1339 , n152 ); 
nand ( n2397 , n2395 , n2396 ); 
nand ( n2398 , n2213 , n2362 ); 
not ( n2399 , n2398 ); 
not ( n2400 , n1261 ); 
or ( n2401 , n2399 , n2400 ); 
not ( n2402 , n149 ); 
or ( n2403 , n1261 , n2402 ); 
nand ( n2404 , n2401 , n2403 ); 
not ( n2405 , n1226 ); 
nand ( n2406 , n2405 , n1229 ); 
not ( n2407 , n2406 ); 
not ( n2408 , n179 ); 
or ( n2409 , n2407 , n2408 ); 
not ( n2410 , n1138 ); 
nand ( n2411 , n127 , n128 , n134 , n142 ); 
nand ( n2412 , n104 , n111 , n115 , n119 ); 
nand ( n2413 , n87 , n92 , n95 , n103 ); 
nor ( n2414 , n2411 , n2412 , n2413 ); 
and ( n2415 , n2410 , n1145 , n2414 ); 
not ( n2416 , n97 ); 
not ( n2417 , n693 ); 
or ( n2418 , n2416 , n2417 ); 
and ( n2419 , n524 , n99 ); 
and ( n2420 , n824 , n98 ); 
nor ( n2421 , n2419 , n2420 ); 
nand ( n2422 , n2418 , n2421 ); 
nor ( n2423 , n2415 , n2422 ); 
or ( n2424 , n2423 , n2406 ); 
nand ( n2425 , n2409 , n2424 ); 
or ( n2426 , n1230 , n1239 ); 
nand ( n2427 , n2426 , n1421 ); 
not ( n2428 , n178 ); 
not ( n2429 , n2406 ); 
or ( n2430 , n2428 , n2429 ); 
or ( n2431 , n2406 , n1115 ); 
nand ( n2432 , n2430 , n2431 ); 
and ( n2433 , n1338 , n2398 ); 
not ( n2434 , n1338 ); 
and ( n2435 , n2434 , n148 ); 
or ( n2436 , n2433 , n2435 ); 
not ( n2437 , n1651 ); 
not ( n2438 , n2062 ); 
or ( n2439 , n2437 , n2438 ); 
nand ( n2440 , n2439 , n2042 ); 
not ( n2441 , n1557 ); 
not ( n2442 , n151 ); 
or ( n2443 , n2441 , n2442 ); 
or ( n2444 , n1262 , n2394 ); 
nand ( n2445 , n2443 , n2444 ); 
not ( n2446 , n56 ); 
not ( n2447 , n1608 ); 
or ( n2448 , n2446 , n2447 ); 
or ( n2449 , n1768 , n1613 ); 
nand ( n2450 , n2448 , n2449 ); 
patch p0 (.t_0(t_0), .g1(n2169), .g2(n1003), .g3(n2207), .g4(n2278), .g5(n2174), .g6(n995), .g7(n1172), .g8(n598), .g9(g238), .g10(n1621), .g11(n2180), .g12(n630), .g13(n323), .g14(n318), .g15(n152), .g16(n604));
endmodule 

