module patch (t_0, t_1, t_2, t_3, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48;
output t_0, t_1, t_2, t_3;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630;

nor ( w1 , g1 , g2 );
nor ( w2 , w1 , g3 );
and ( w3 , w2 , w6138 );
and ( w4 , w51 , g5 );
nor ( w5 , g5 , g6 );
nor ( w6 , w4 , w5 );
nor ( w7 , w6 , g7 );
nor ( w8 , g7 , g5 );
and ( w9 , g6 , w8 );
nor ( w10 , g4 , g3 );
and ( w11 , w3175 , w10 );
and ( w12 , w11 , g7 );
nor ( w13 , w12 , w9 );
and ( w14 , w11 , g5 );
and ( w15 , w13 , w6148 );
not ( w16 , w9 );
and ( w17 , w16 , w15 );
and ( w18 , g8 , g9 );
and ( w19 , g10 , g11 );
nor ( w20 , g12 , g13 );
and ( w21 , g14 , g15 );
nor ( w22 , w21 , g16 );
and ( w23 , g14 , g16 );
and ( w24 , w23 , g15 );
nor ( w25 , w24 , g17 );
nor ( w26 , w22 , w25 );
nor ( w27 , w26 , g18 );
and ( w28 , w26 , g18 );
nor ( w29 , w28 , g19 );
nor ( w30 , w27 , w29 );
nor ( w31 , g20 , g21 );
and ( w32 , w30 , w7485 );
and ( w33 , g22 , g23 );
nor ( w34 , w32 , w33 );
and ( w35 , g20 , g21 );
and ( w36 , w34 , w8363 );
nor ( w37 , g22 , g23 );
nor ( w38 , w36 , w37 );
and ( w39 , g24 , g25 );
nor ( w40 , w38 , w39 );
nor ( w41 , g24 , g25 );
nor ( w42 , w40 , w41 );
nor ( w43 , g26 , g27 );
and ( w44 , w42 , w12144 );
and ( w45 , g26 , g27 );
nor ( w46 , w44 , w45 );
and ( w47 , w46 , w12919 );
nor ( w48 , g8 , g9 );
and ( w49 , w48 , w12919 );
nor ( w50 , w49 , w20 );
not ( w51 , w3 );
and ( w52 , w51 , g7 );
nor ( w53 , w7 , w52 );
nor ( w54 , w50 , w53 );
nor ( w55 , w47 , w54 );
and ( w56 , g17 , g16 );
not ( w57 , w56 );
and ( w58 , w57 , g16 );
not ( w59 , w58 );
and ( w60 , w59 , g17 );
not ( w61 , w60 );
and ( w62 , w61 , g17 );
nor ( w63 , w62 , w35 );
and ( w64 , w63 , w12424 );
nor ( w65 , w1 , g2 );
and ( w66 , w65 , w2636 );
and ( w67 , w2562 , w10 );
nor ( w68 , w67 , g3 );
and ( w69 , w68 , w6138 );
nor ( w70 , w66 , g3 );
and ( w71 , w70 , w6138 );
nor ( w72 , w71 , g3 );
and ( w73 , w72 , w6138 );
nor ( w74 , w69 , w73 );
nor ( w75 , w5 , w52 );
and ( w76 , w75 , w11092 );
nor ( w77 , w76 , w53 );
and ( w78 , w74 , w77 );
and ( w79 , w78 , w12612 );
and ( w80 , w64 , w79 );
nor ( w81 , w37 , w80 );
nor ( w82 , w81 , w33 );
and ( w83 , w82 , w12144 );
and ( w84 , w83 , w7803 );
and ( w85 , w84 , w79 );
nor ( w86 , w41 , w85 );
and ( w87 , w86 , w12144 );
nor ( w88 , w87 , w45 );
nor ( w89 , w20 , w88 );
and ( w90 , w89 , w12142 );
not ( w91 , w90 );
and ( w92 , w91 , w79 );
and ( w93 , w92 , w12612 );
and ( w94 , w257 , w93 );
and ( w95 , w12921 , g9 );
and ( w96 , w95 , g8 );
not ( w97 , w96 );
and ( w98 , w97 , g8 );
and ( w99 , w98 , g9 );
not ( w100 , w99 );
and ( w101 , w100 , w18 );
and ( w102 , w101 , w12612 );
nor ( w103 , w94 , w102 );
nor ( w104 , w103 , w18 );
and ( w105 , g12 , g13 );
and ( w106 , w104 , w11166 );
and ( w107 , w106 , w79 );
and ( w108 , w107 , w12612 );
and ( w109 , w1573 , w108 );
and ( w110 , w109 , w48 );
and ( w111 , w11166 , w15 );
not ( w112 , w110 );
and ( w113 , w112 , w111 );
and ( w114 , w113 , w203 );
and ( w115 , w114 , w17 );
and ( w116 , w115 , w15 );
not ( w117 , w116 );
and ( w118 , w117 , w79 );
and ( w119 , w118 , w48 );
and ( w120 , w119 , w79 );
and ( w121 , w118 , w120 );
not ( w122 , w121 );
and ( w123 , w122 , w48 );
and ( w124 , w39 , w17 );
and ( w125 , w12142 , w17 );
and ( w126 , w124 , w125 );
nor ( w127 , w126 , w43 );
not ( w128 , w127 );
and ( w129 , w128 , w17 );
and ( w130 , w12144 , w17 );
and ( w131 , w129 , w130 );
and ( w132 , w131 , w12921 );
and ( w133 , w132 , w17 );
and ( w134 , w12057 , g29 );
not ( w135 , w134 );
and ( w136 , w135 , g29 );
and ( w137 , w136 , w17 );
nor ( w138 , w133 , w137 );
and ( w139 , w138 , g30 );
not ( w140 , w139 );
and ( w141 , w140 , g30 );
not ( w142 , w141 );
and ( w143 , w142 , g31 );
not ( w144 , w143 );
and ( w145 , w144 , g31 );
and ( w146 , w33 , w7803 );
and ( w147 , w39 , w7803 );
not ( w148 , w147 );
and ( w149 , w148 , w37 );
and ( w150 , w149 , w12117 );
and ( w151 , w21 , g17 );
and ( w152 , w21 , g16 );
nor ( w153 , w151 , w152 );
and ( w154 , w7485 , g17 );
and ( w155 , w154 , g16 );
and ( w156 , w155 , g18 );
and ( w157 , w156 , g17 );
nor ( w158 , w157 , w39 );
and ( w159 , w158 , w11347 );
and ( w160 , w153 , w159 );
and ( w161 , w160 , w9197 );
not ( w162 , w161 );
and ( w163 , w162 , g18 );
and ( w164 , w261 , g17 );
nor ( w165 , w164 , w152 );
not ( w166 , w165 );
and ( w167 , w166 , g19 );
nor ( w168 , w163 , w167 );
nor ( w169 , w168 , w31 );
nor ( w170 , w169 , w35 );
and ( w171 , w170 , w11140 );
and ( w172 , w11347 , w171 );
nor ( w173 , w172 , w41 );
nor ( w174 , w173 , w45 );
nor ( w175 , w150 , w174 );
and ( w176 , w175 , w12921 );
and ( w177 , w176 , w12144 );
and ( w178 , w177 , w12142 );
and ( w179 , w178 , w12612 );
not ( w180 , w179 );
and ( w181 , w146 , w180 );
and ( w182 , w181 , w12144 );
and ( w183 , w182 , w17 );
nor ( w184 , w183 , w45 );
nor ( w185 , w184 , w179 );
and ( w186 , w185 , w17 );
nor ( w187 , w186 , w45 );
nor ( w188 , w187 , w179 );
and ( w189 , w188 , w17 );
nor ( w190 , w189 , w45 );
nor ( w191 , w40 , w43 );
nor ( w192 , w191 , w18 );
nor ( w193 , w192 , w41 );
nor ( w194 , w45 , w18 );
nor ( w195 , w48 , w20 );
nor ( w196 , w195 , w53 );
nor ( w197 , w194 , w196 );
nor ( w198 , w193 , w197 );
nor ( w199 , w198 , w196 );
not ( w200 , w199 );
and ( w201 , w190 , w200 );
nor ( w202 , w201 , w179 );
not ( w203 , w102 );
and ( w204 , w202 , w203 );
and ( w205 , w204 , w17 );
and ( w206 , w7402 , g7 );
nor ( w207 , w5 , g6 );
and ( w208 , w207 , w11092 );
and ( w209 , g6 , w77 );
nor ( w210 , w209 , w52 );
and ( w211 , w210 , w11092 );
and ( w212 , w12934 , w5 );
and ( w213 , w211 , w7419 );
nor ( w214 , w213 , g5 );
nor ( w215 , g5 , w214 );
nor ( w216 , w215 , w53 );
and ( w217 , w7402 , w216 );
and ( w218 , g6 , w11092 );
and ( w219 , w12934 , w218 );
not ( w220 , w219 );
and ( w221 , w220 , w1 );
and ( w222 , w10 , g7 );
nor ( w223 , w222 , w219 );
and ( w224 , w10 , g5 );
and ( w225 , w223 , w7415 );
nor ( w226 , w221 , w225 );
nor ( w227 , w217 , w226 );
nor ( w228 , w208 , w227 );
and ( w229 , w228 , w12934 );
nor ( w230 , w206 , w229 );
nor ( w231 , w205 , w230 );
and ( w232 , w231 , w12612 );
not ( w233 , w145 );
and ( w234 , w233 , w232 );
and ( w235 , w11140 , w41 );
and ( w236 , w33 , w17 );
and ( w237 , w12424 , w17 );
nor ( w238 , w236 , w237 );
nor ( w239 , w33 , w35 );
nor ( w240 , w238 , w239 );
nor ( w241 , w240 , w39 );
not ( w242 , w241 );
and ( w243 , w242 , w17 );
and ( w244 , w12144 , w243 );
not ( w245 , w235 );
and ( w246 , w245 , w244 );
and ( w247 , w234 , w368 );
and ( w248 , w247 , w12117 );
and ( w249 , w38 , w12144 );
and ( w250 , w249 , w7803 );
not ( w251 , w250 );
and ( w252 , w248 , w251 );
nor ( w253 , w48 , w252 );
and ( w254 , w253 , w125 );
and ( w255 , g28 , g29 );
nor ( w256 , w254 , w255 );
not ( w257 , w55 );
and ( w258 , w256 , w257 );
not ( w259 , w25 );
and ( w260 , w259 , w17 );
not ( w261 , w22 );
and ( w262 , w261 , w260 );
and ( w263 , w262 , w17 );
and ( w264 , w263 , w15 );
and ( w265 , w264 , w17 );
and ( w266 , w265 , w15 );
and ( w267 , w260 , w266 );
and ( w268 , w267 , w17 );
and ( w269 , w268 , w15 );
and ( w270 , w21 , w269 );
nor ( w271 , w270 , w56 );
and ( w272 , g18 , g19 );
and ( w273 , w271 , w12085 );
nor ( w274 , g18 , g19 );
and ( w275 , w3811 , w17 );
not ( w276 , w273 );
and ( w277 , w276 , w275 );
nor ( w278 , w277 , w171 );
not ( w279 , w278 );
and ( w280 , w279 , w17 );
and ( w281 , w280 , w8363 );
and ( w282 , w281 , w11347 );
nor ( w283 , w41 , w282 );
not ( w284 , w283 );
and ( w285 , w284 , w237 );
nor ( w286 , w285 , w124 );
and ( w287 , w286 , w368 );
and ( w288 , w287 , w12424 );
and ( w289 , w288 , w12117 );
and ( w290 , w39 , w1935 );
not ( w291 , w290 );
and ( w292 , w291 , w125 );
not ( w293 , w292 );
and ( w294 , w293 , w179 );
not ( w295 , w294 );
and ( w296 , w295 , w17 );
not ( w297 , w289 );
and ( w298 , w297 , w296 );
and ( w299 , w298 , w130 );
nor ( w300 , w43 , w299 );
not ( w301 , w300 );
and ( w302 , w301 , w17 );
nor ( w303 , w302 , w230 );
and ( w304 , w303 , w12612 );
nor ( w305 , w258 , w304 );
nor ( w306 , w20 , w305 );
and ( w307 , w306 , w8848 );
nor ( w308 , g32 , g33 );
and ( w309 , w12532 , w17 );
and ( w310 , g30 , g31 );
and ( w311 , w310 , w17 );
and ( w312 , g32 , g33 );
and ( w313 , w308 , w12037 );
and ( w314 , w311 , w313 );
and ( w315 , w314 , w308 );
not ( w316 , w315 );
and ( w317 , w316 , w310 );
nor ( w318 , w317 , w312 );
and ( w319 , w312 , w17 );
nor ( w320 , w318 , w319 );
and ( w321 , w12080 , w320 );
nor ( w322 , w313 , w309 );
not ( w323 , w322 );
and ( w324 , w323 , w17 );
and ( w325 , w324 , w15 );
not ( w326 , w321 );
and ( w327 , w326 , w325 );
and ( w328 , w327 , w17 );
nor ( w329 , w328 , w230 );
and ( w330 , w329 , w79 );
and ( w331 , w330 , w12612 );
and ( w332 , w1064 , w331 );
nor ( w333 , w17 , w230 );
and ( w334 , w333 , w12612 );
nor ( w335 , w332 , w334 );
and ( w336 , w335 , g30 );
and ( w337 , w336 , g31 );
not ( w338 , w337 );
and ( w339 , w338 , w310 );
and ( w340 , g34 , g35 );
not ( w341 , w340 );
and ( w342 , w341 , g34 );
not ( w343 , w342 );
and ( w344 , w343 , g34 );
not ( w345 , w344 );
and ( w346 , w345 , g35 );
not ( w347 , w346 );
and ( w348 , w347 , g35 );
and ( w349 , w12381 , g34 );
not ( w350 , w349 );
and ( w351 , g34 , w350 );
not ( w352 , w348 );
and ( w353 , w352 , w351 );
and ( w354 , w353 , w12612 );
not ( w355 , w230 );
and ( w356 , w354 , w355 );
and ( w357 , w356 , w12612 );
nor ( w358 , w339 , w357 );
not ( w359 , w304 );
and ( w360 , w358 , w359 );
nor ( w361 , w255 , w360 );
not ( w362 , w361 );
and ( w363 , w362 , w325 );
nor ( w364 , w282 , w37 );
and ( w365 , w7803 , w364 );
not ( w366 , w124 );
and ( w367 , w365 , w366 );
not ( w368 , w246 );
and ( w369 , w367 , w368 );
and ( w370 , w12117 , w369 );
nor ( w371 , w370 , w48 );
nor ( w372 , w371 , w43 );
and ( w373 , w372 , w12142 );
and ( w374 , w216 , w79 );
nor ( w375 , w374 , w226 );
nor ( w376 , w375 , w255 );
nor ( w377 , g28 , g29 );
and ( w378 , w255 , w12498 );
not ( w379 , w378 );
and ( w380 , w379 , w17 );
and ( w381 , w555 , w255 );
not ( w382 , w381 );
and ( w383 , w382 , w17 );
nor ( w384 , g30 , g31 );
nor ( w385 , w383 , w384 );
nor ( w386 , w375 , w310 );
and ( w387 , w386 , w384 );
not ( w388 , w387 );
and ( w389 , w388 , w15 );
not ( w390 , w385 );
and ( w391 , w390 , w389 );
not ( w392 , w391 );
and ( w393 , w392 , w255 );
and ( w394 , w393 , w216 );
and ( w395 , w394 , w79 );
and ( w396 , w395 , w12612 );
nor ( w397 , w376 , w396 );
nor ( w398 , w19 , w397 );
not ( w399 , w15 );
and ( w400 , w377 , w399 );
and ( w401 , w19 , w400 );
nor ( w402 , w401 , g12 );
and ( w403 , w402 , w111 );
and ( w404 , w403 , w20 );
and ( w405 , w404 , w11797 );
and ( w406 , w405 , w20 );
and ( w407 , w12379 , g35 );
nor ( w408 , w407 , w349 );
and ( w409 , w408 , w79 );
and ( w410 , w408 , w79 );
nor ( w411 , w409 , w410 );
not ( w412 , w400 );
and ( w413 , w412 , w411 );
nor ( w414 , w48 , w17 );
nor ( w415 , w35 , w236 );
not ( w416 , w415 );
and ( w417 , w416 , w237 );
and ( w418 , w39 , w15 );
nor ( w419 , w417 , w418 );
not ( w420 , w419 );
and ( w421 , w420 , w17 );
and ( w422 , w421 , w15 );
nor ( w423 , w37 , w422 );
not ( w424 , w423 );
and ( w425 , w424 , w243 );
and ( w426 , w425 , w11140 );
nor ( w427 , w426 , w418 );
nor ( w428 , g16 , g17 );
and ( w429 , w11132 , w21 );
nor ( w430 , w429 , w56 );
and ( w431 , w430 , w12085 );
and ( w432 , w272 , w15 );
and ( w433 , w432 , g19 );
and ( w434 , w7485 , w432 );
nor ( w435 , w434 , w35 );
not ( w436 , w435 );
and ( w437 , w436 , w17 );
and ( w438 , w437 , w15 );
and ( w439 , w433 , w438 );
and ( w440 , w439 , w11347 );
and ( w441 , w440 , w17 );
and ( w442 , w441 , w15 );
nor ( w443 , w266 , w442 );
not ( w444 , w431 );
and ( w445 , w444 , w443 );
and ( w446 , w445 , w3811 );
nor ( w447 , w446 , w35 );
and ( w448 , w7485 , w15 );
and ( w449 , w447 , w448 );
and ( w450 , w449 , w237 );
nor ( w451 , w450 , w31 );
and ( w452 , w451 , w12424 );
nor ( w453 , w452 , w33 );
and ( w454 , w453 , w17 );
and ( w455 , w454 , w15 );
not ( w456 , w226 );
and ( w457 , w455 , w456 );
and ( w458 , w457 , w11140 );
not ( w459 , w458 );
and ( w460 , w459 , w427 );
not ( w461 , w418 );
and ( w462 , w460 , w461 );
nor ( w463 , w462 , w226 );
not ( w464 , w463 );
and ( w465 , w427 , w464 );
and ( w466 , w7803 , w15 );
and ( w467 , w961 , w466 );
nor ( w468 , w467 , w41 );
nor ( w469 , w468 , w45 );
and ( w470 , w45 , w15 );
nor ( w471 , w469 , w470 );
not ( w472 , w471 );
and ( w473 , w472 , w130 );
nor ( w474 , w473 , w43 );
not ( w475 , w474 );
and ( w476 , w475 , w15 );
nor ( w477 , w476 , w53 );
nor ( w478 , w414 , w477 );
and ( w479 , w478 , w12919 );
and ( w480 , w18 , w15 );
nor ( w481 , w479 , w480 );
not ( w482 , w481 );
and ( w483 , w482 , w15 );
and ( w484 , w413 , w483 );
nor ( w485 , g10 , g11 );
nor ( w486 , w485 , w226 );
and ( w487 , w484 , w486 );
and ( w488 , w487 , w19 );
nor ( w489 , w216 , w226 );
and ( w490 , w20 , w1231 );
nor ( w491 , w375 , w489 );
and ( w492 , w491 , w216 );
and ( w493 , w492 , w79 );
nor ( w494 , w493 , w226 );
and ( w495 , w1231 , w79 );
nor ( w496 , w495 , w226 );
nor ( w497 , w494 , w496 );
and ( w498 , w497 , w1231 );
and ( w499 , w498 , w216 );
and ( w500 , w499 , w79 );
nor ( w501 , w500 , w226 );
nor ( w502 , w79 , w226 );
nor ( w503 , w501 , w502 );
and ( w504 , w503 , w1231 );
and ( w505 , w504 , w216 );
and ( w506 , w505 , w79 );
nor ( w507 , w506 , w226 );
not ( w508 , w507 );
and ( w509 , w508 , w216 );
and ( w510 , w509 , w79 );
nor ( w511 , w510 , w226 );
not ( w512 , w511 );
and ( w513 , w512 , w216 );
and ( w514 , w513 , w79 );
nor ( w515 , w514 , w226 );
nor ( w516 , w515 , w501 );
and ( w517 , w516 , w1231 );
and ( w518 , w517 , w12144 );
not ( w519 , w518 );
and ( w520 , w519 , w111 );
and ( w521 , w520 , w12919 );
and ( w522 , w8640 , w15 );
and ( w523 , w522 , w480 );
nor ( w524 , w521 , w523 );
and ( w525 , w524 , w1055 );
not ( w526 , w525 );
and ( w527 , w526 , w15 );
not ( w528 , w527 );
and ( w529 , w528 , w216 );
and ( w530 , w529 , w79 );
and ( w531 , w530 , w12612 );
nor ( w532 , w490 , w531 );
nor ( w533 , w532 , w375 );
and ( w534 , w533 , w12612 );
nor ( w535 , w534 , w20 );
nor ( w536 , w501 , w375 );
not ( w537 , w535 );
and ( w538 , w537 , w536 );
not ( w539 , w538 );
and ( w540 , w539 , w15 );
not ( w541 , w540 );
and ( w542 , w541 , w216 );
and ( w543 , w542 , w79 );
and ( w544 , w543 , w12612 );
and ( w545 , w1055 , w544 );
and ( w546 , w545 , w12612 );
and ( w547 , w538 , w546 );
not ( w548 , w547 );
and ( w549 , w548 , w15 );
not ( w550 , w549 );
and ( w551 , w550 , w216 );
and ( w552 , w551 , w79 );
and ( w553 , w552 , w12612 );
and ( w554 , w553 , w12080 );
not ( w555 , w380 );
and ( w556 , w536 , w555 );
and ( w557 , w556 , w485 );
and ( w558 , w557 , w12142 );
and ( w559 , w558 , w1452 );
and ( w560 , w12142 , w559 );
nor ( w561 , w560 , w20 );
nor ( w562 , w561 , w489 );
and ( w563 , w562 , w216 );
and ( w564 , w563 , w79 );
and ( w565 , w564 , w12612 );
and ( w566 , w565 , w11166 );
and ( w567 , w566 , w216 );
and ( w568 , w567 , w12612 );
and ( w569 , w568 , w12717 );
and ( w570 , w569 , w384 );
and ( w571 , w570 , w11166 );
not ( w572 , w571 );
and ( w573 , w572 , w15 );
not ( w574 , w573 );
and ( w575 , w574 , w79 );
and ( w576 , w575 , w12612 );
nor ( w577 , w385 , w576 );
not ( w578 , w577 );
and ( w579 , w578 , w255 );
and ( w580 , w579 , w11166 );
and ( w581 , w580 , w79 );
and ( w582 , w581 , w12612 );
nor ( w583 , w582 , w20 );
nor ( w584 , w583 , w489 );
and ( w585 , w584 , w12612 );
nor ( w586 , w554 , w585 );
and ( w587 , w554 , w377 );
and ( w588 , w12142 , w587 );
not ( w589 , w588 );
and ( w590 , w589 , w483 );
and ( w591 , w590 , w12919 );
not ( w592 , w591 );
and ( w593 , w592 , w485 );
and ( w594 , w593 , w1452 );
not ( w595 , w594 );
and ( w596 , w595 , w111 );
nor ( w597 , w596 , w105 );
nor ( w598 , w111 , w486 );
not ( w599 , w598 );
and ( w600 , w599 , w15 );
not ( w601 , w597 );
and ( w602 , w601 , w600 );
and ( w603 , w411 , w483 );
and ( w604 , w603 , w125 );
nor ( w605 , w604 , w48 );
not ( w606 , w605 );
and ( w607 , w606 , w111 );
and ( w608 , w15 , w411 );
and ( w609 , w608 , w600 );
and ( w610 , w609 , w105 );
and ( w611 , w610 , w8640 );
and ( w612 , w611 , w522 );
and ( w613 , w612 , w105 );
and ( w614 , w613 , w8848 );
and ( w615 , w614 , w12921 );
and ( w616 , w615 , w12037 );
not ( w617 , w408 );
and ( w618 , w617 , g32 );
and ( w619 , w618 , g33 );
nor ( w620 , w619 , w308 );
and ( w621 , w620 , w79 );
nor ( w622 , w408 , w621 );
and ( w623 , w622 , w15 );
nor ( w624 , g34 , g35 );
nor ( w625 , w624 , g35 );
nor ( w626 , w625 , w407 );
not ( w627 , w407 );
and ( w628 , w627 , g35 );
nor ( w629 , w628 , w624 );
nor ( w630 , w407 , w629 );
not ( w631 , w630 );
and ( w632 , w631 , w216 );
and ( w633 , w626 , w699 );
and ( w634 , w349 , w216 );
nor ( w635 , w634 , w632 );
and ( w636 , w377 , w635 );
and ( w637 , w636 , w13333 );
not ( w638 , w637 );
and ( w639 , w638 , w377 );
not ( w640 , w633 );
and ( w641 , w640 , w216 );
nor ( w642 , w639 , w641 );
and ( w643 , w642 , w15 );
and ( w644 , w633 , w643 );
and ( w645 , w644 , w19 );
nor ( w646 , w384 , g30 );
nor ( w647 , w646 , g31 );
nor ( w648 , w647 , g31 );
nor ( w649 , w383 , w648 );
and ( w650 , w649 , w11852 );
and ( w651 , w12717 , w384 );
not ( w652 , w651 );
and ( w653 , w652 , w15 );
not ( w654 , w650 );
and ( w655 , w654 , w653 );
not ( w656 , w655 );
and ( w657 , w656 , w255 );
nor ( w658 , w657 , w19 );
not ( w659 , w658 );
and ( w660 , w659 , w79 );
and ( w661 , w660 , w12612 );
nor ( w662 , w376 , w661 );
not ( w663 , w662 );
and ( w664 , w663 , w216 );
and ( w665 , w664 , w79 );
and ( w666 , w665 , w12612 );
not ( w667 , w645 );
and ( w668 , w667 , w666 );
nor ( w669 , w668 , g12 );
and ( w670 , w669 , w111 );
not ( w671 , w670 );
and ( w672 , w671 , w93 );
nor ( w673 , w672 , g13 );
and ( w674 , w673 , w20 );
and ( w675 , w678 , w216 );
nor ( w676 , w675 , w310 );
nor ( w677 , w310 , w255 );
not ( w678 , w626 );
and ( w679 , w678 , w216 );
nor ( w680 , w677 , w679 );
and ( w681 , w680 , w11852 );
nor ( w682 , w681 , w648 );
and ( w683 , w682 , w79 );
not ( w684 , w676 );
and ( w685 , w684 , w683 );
nor ( w686 , w632 , w685 );
and ( w687 , w626 , w769 );
not ( w688 , w675 );
and ( w689 , w687 , w688 );
not ( w690 , w689 );
and ( w691 , w690 , w216 );
not ( w692 , w691 );
and ( w693 , w687 , w692 );
not ( w694 , w693 );
and ( w695 , w694 , w216 );
nor ( w696 , w695 , w632 );
not ( w697 , w685 );
and ( w698 , w697 , w696 );
not ( w699 , w632 );
and ( w700 , w698 , w699 );
and ( w701 , w696 , w105 );
not ( w702 , w696 );
and ( w703 , w377 , w702 );
not ( w704 , w703 );
and ( w705 , w704 , w700 );
and ( w706 , w705 , w12921 );
and ( w707 , w706 , w105 );
not ( w708 , w707 );
and ( w709 , w708 , g13 );
not ( w710 , w709 );
and ( w711 , w710 , g13 );
and ( w712 , w491 , w8848 );
and ( w713 , w712 , w20 );
and ( w714 , w713 , w79 );
and ( w715 , w714 , w12612 );
and ( w716 , w12717 , w715 );
and ( w717 , w716 , w1055 );
and ( w718 , w717 , w1231 );
and ( w719 , w718 , w20 );
and ( w720 , w719 , w12080 );
and ( w721 , w720 , w8848 );
nor ( w722 , w477 , w18 );
nor ( w723 , w722 , w480 );
not ( w724 , w723 );
and ( w725 , w724 , w377 );
and ( w726 , w725 , w13333 );
and ( w727 , w726 , w15 );
and ( w728 , w727 , w8848 );
and ( w729 , w467 , w12117 );
nor ( w730 , w729 , w470 );
not ( w731 , w730 );
and ( w732 , w731 , w130 );
nor ( w733 , w732 , w43 );
and ( w734 , w733 , w179 );
nor ( w735 , w734 , w102 );
and ( w736 , w735 , w12919 );
nor ( w737 , w736 , w480 );
nor ( w738 , w737 , w351 );
nor ( w739 , w738 , g35 );
not ( w740 , w739 );
and ( w741 , w740 , w377 );
and ( w742 , w748 , w377 );
not ( w743 , w354 );
and ( w744 , w742 , w743 );
and ( w745 , w744 , w15 );
nor ( w746 , w745 , w53 );
and ( w747 , w744 , w763 );
not ( w748 , w737 );
and ( w749 , w748 , w15 );
nor ( w750 , w749 , w53 );
nor ( w751 , w737 , w750 );
and ( w752 , w751 , w15 );
nor ( w753 , w752 , w53 );
not ( w754 , w753 );
and ( w755 , w747 , w754 );
and ( w756 , w755 , w377 );
and ( w757 , w756 , w13333 );
and ( w758 , w757 , w15 );
nor ( w759 , w758 , w53 );
not ( w760 , w759 );
and ( w761 , w741 , w760 );
and ( w762 , w761 , w763 );
not ( w763 , w746 );
and ( w764 , w742 , w763 );
and ( w765 , w764 , w15 );
nor ( w766 , w765 , w53 );
not ( w767 , w766 );
and ( w768 , w762 , w767 );
not ( w769 , w634 );
and ( w770 , w768 , w769 );
not ( w771 , w770 );
and ( w772 , w771 , w377 );
nor ( w773 , w772 , w685 );
not ( w774 , w773 );
and ( w775 , w19 , w774 );
not ( w776 , w775 );
and ( w777 , w776 , w15 );
not ( w778 , w777 );
and ( w779 , w778 , w79 );
and ( w780 , w779 , w12612 );
not ( w781 , w780 );
and ( w782 , w781 , w19 );
and ( w783 , w782 , w15 );
not ( w784 , w783 );
and ( w785 , w784 , w79 );
not ( w786 , w728 );
and ( w787 , w786 , w785 );
and ( w788 , w715 , w1055 );
nor ( w789 , w377 , w255 );
and ( w790 , w5536 , g30 );
not ( w791 , w790 );
and ( w792 , w791 , g30 );
not ( w793 , w792 );
and ( w794 , w793 , g31 );
not ( w795 , w794 );
and ( w796 , w795 , g31 );
not ( w797 , w796 );
and ( w798 , w797 , w79 );
and ( w799 , w788 , w798 );
and ( w800 , w799 , w1055 );
and ( w801 , w800 , w1573 );
nor ( w802 , w801 , w179 );
not ( w803 , w802 );
and ( w804 , w20 , w803 );
not ( w805 , w804 );
and ( w806 , w805 , w377 );
nor ( w807 , w19 , w806 );
not ( w808 , w807 );
and ( w809 , w808 , w377 );
nor ( w810 , w809 , g29 );
not ( w811 , w810 );
and ( w812 , w811 , w377 );
and ( w813 , w812 , w13333 );
and ( w814 , w813 , w111 );
and ( w815 , w814 , w125 );
nor ( w816 , w815 , w48 );
not ( w817 , w816 );
and ( w818 , w817 , w15 );
not ( w819 , w818 );
and ( w820 , w819 , w216 );
and ( w821 , w820 , w79 );
and ( w822 , w821 , w12612 );
nor ( w823 , w787 , w822 );
and ( w824 , w377 , w19 );
nor ( w825 , w824 , w375 );
and ( w826 , w825 , w312 );
and ( w827 , w825 , w1064 );
and ( w828 , w827 , w13211 );
not ( w829 , w828 );
and ( w830 , w829 , w377 );
and ( w831 , w830 , w13333 );
and ( w832 , w831 , w15 );
not ( w833 , w826 );
and ( w834 , w833 , w832 );
nor ( w835 , w834 , w489 );
and ( w836 , w835 , w20 );
not ( w837 , w468 );
and ( w838 , w837 , w130 );
nor ( w839 , w838 , w43 );
not ( w840 , w839 );
and ( w841 , w840 , w377 );
and ( w842 , w841 , w12919 );
nor ( w843 , w842 , w480 );
not ( w844 , w843 );
and ( w845 , w844 , w377 );
nor ( w846 , w845 , w45 );
and ( w847 , w377 , w522 );
nor ( w848 , w847 , w375 );
and ( w849 , w848 , g30 );
and ( w850 , w849 , w13206 );
and ( w851 , w848 , w12199 );
and ( w852 , w851 , g31 );
not ( w853 , w852 );
and ( w854 , w853 , w15 );
not ( w855 , w850 );
and ( w856 , w855 , w854 );
not ( w857 , w856 );
and ( w858 , w857 , g26 );
not ( w859 , w858 );
and ( w860 , w859 , g26 );
not ( w861 , w860 );
and ( w862 , w861 , g27 );
not ( w863 , w862 );
and ( w864 , w863 , w470 );
and ( w865 , w864 , g27 );
nor ( w866 , w865 , w43 );
and ( w867 , w866 , w45 );
not ( w868 , w867 );
and ( w869 , w868 , w15 );
not ( w870 , w869 );
and ( w871 , w870 , w216 );
and ( w872 , w871 , w79 );
and ( w873 , w872 , w12612 );
nor ( w874 , w846 , w873 );
nor ( w875 , w19 , w874 );
and ( w876 , w470 , g27 );
and ( w877 , w626 , w12498 );
and ( w878 , w377 , w105 );
nor ( w879 , w878 , w125 );
and ( w880 , w847 , w15 );
and ( w881 , w880 , w522 );
and ( w882 , w881 , w377 );
and ( w883 , w882 , w13333 );
and ( w884 , w883 , w15 );
not ( w885 , w879 );
and ( w886 , w885 , w884 );
and ( w887 , w886 , w8848 );
and ( w888 , w887 , w522 );
and ( w889 , w888 , w17 );
and ( w890 , w889 , w15 );
nor ( w891 , w877 , w890 );
and ( w892 , w891 , w8848 );
and ( w893 , w377 , w414 );
and ( w894 , w19 , w893 );
not ( w895 , w894 );
and ( w896 , w895 , w17 );
and ( w897 , w896 , w15 );
not ( w898 , w892 );
and ( w899 , w898 , w897 );
and ( w900 , w961 , w899 );
not ( w901 , w629 );
and ( w902 , w900 , w901 );
and ( w903 , w120 , w11166 );
and ( w904 , w903 , w8848 );
and ( w905 , w904 , w79 );
nor ( w906 , w905 , w226 );
and ( w907 , w902 , w906 );
and ( w908 , w907 , w466 );
nor ( w909 , w908 , w41 );
not ( w910 , w909 );
and ( w911 , w910 , w130 );
nor ( w912 , w911 , w43 );
nor ( w913 , w19 , w377 );
and ( w914 , w19 , w12498 );
not ( w915 , w914 );
and ( w916 , w915 , w17 );
and ( w917 , w916 , w15 );
not ( w918 , w913 );
and ( w919 , w918 , w917 );
not ( w920 , w919 );
and ( w921 , w920 , w377 );
nor ( w922 , w921 , w629 );
and ( w923 , w922 , w17 );
and ( w924 , w923 , w15 );
not ( w925 , w912 );
and ( w926 , w925 , w924 );
and ( w927 , w926 , w12117 );
nor ( w928 , w927 , w255 );
nor ( w929 , w928 , w485 );
and ( w930 , w929 , w522 );
and ( w931 , w930 , w12919 );
and ( w932 , w931 , w12080 );
and ( w933 , w932 , w17 );
and ( w934 , w933 , w15 );
not ( w935 , w934 );
and ( w936 , w935 , w216 );
and ( w937 , w936 , w79 );
nor ( w938 , w937 , w226 );
nor ( w939 , w876 , w938 );
not ( w940 , w480 );
and ( w941 , w939 , w940 );
and ( w942 , w941 , w13206 );
nor ( w943 , w942 , w746 );
and ( w944 , w943 , w377 );
not ( w945 , w944 );
and ( w946 , w19 , w945 );
and ( w947 , w946 , w312 );
and ( w948 , w12921 , w947 );
and ( w949 , w948 , w13333 );
not ( w950 , w949 );
and ( w951 , w950 , w377 );
and ( w952 , w951 , w13333 );
and ( w953 , w952 , w15 );
not ( w954 , w953 );
and ( w955 , w954 , w79 );
and ( w956 , w955 , w12612 );
nor ( w957 , w875 , w956 );
and ( w958 , w957 , w924 );
not ( w959 , w958 );
and ( w960 , w959 , w312 );
not ( w961 , w465 );
and ( w962 , w961 , w377 );
and ( w963 , w962 , w466 );
nor ( w964 , w963 , w41 );
not ( w965 , w964 );
and ( w966 , w965 , w130 );
nor ( w967 , w966 , w43 );
nor ( w968 , w967 , w18 );
nor ( w969 , w968 , w480 );
not ( w970 , w969 );
and ( w971 , w970 , w377 );
nor ( w972 , w971 , w45 );
nor ( w973 , w972 , w873 );
nor ( w974 , w973 , w309 );
and ( w975 , w974 , w13211 );
and ( w976 , w8848 , w975 );
nor ( w977 , w976 , w780 );
and ( w978 , w977 , w377 );
and ( w979 , w978 , w13333 );
and ( w980 , w979 , w15 );
not ( w981 , w980 );
and ( w982 , w981 , w79 );
and ( w983 , w982 , w12612 );
nor ( w984 , w960 , w983 );
nor ( w985 , w20 , w984 );
not ( w986 , w985 );
and ( w987 , w986 , w377 );
and ( w988 , w987 , w13333 );
nor ( w989 , w988 , w48 );
not ( w990 , w989 );
and ( w991 , w990 , w125 );
nor ( w992 , w991 , w48 );
not ( w993 , w992 );
and ( w994 , w993 , w15 );
not ( w995 , w994 );
and ( w996 , w995 , w216 );
and ( w997 , w996 , w79 );
and ( w998 , w997 , w12612 );
nor ( w999 , w836 , w998 );
and ( w1000 , w999 , w377 );
and ( w1001 , w1000 , w13333 );
and ( w1002 , w1001 , w15 );
not ( w1003 , w1002 );
and ( w1004 , w1003 , w79 );
and ( w1005 , w1004 , w12612 );
not ( w1006 , w1005 );
and ( w1007 , w823 , w1006 );
nor ( w1008 , w1007 , w255 );
not ( w1009 , w1008 );
and ( w1010 , w377 , w1009 );
and ( w1011 , w1010 , w13333 );
not ( w1012 , w1011 );
and ( w1013 , w1012 , w377 );
nor ( w1014 , w629 , w634 );
not ( w1015 , w1014 );
and ( w1016 , w1015 , w216 );
nor ( w1017 , w1016 , w715 );
not ( w1018 , w1017 );
and ( w1019 , w1018 , w384 );
and ( w1020 , w1231 , w310 );
and ( w1021 , w1020 , w1055 );
and ( w1022 , w1021 , w1231 );
and ( w1023 , w1022 , w20 );
and ( w1024 , w1023 , g32 );
not ( w1025 , w502 );
and ( w1026 , w1024 , w1025 );
and ( w1027 , w1026 , g33 );
and ( w1028 , w1027 , w8848 );
and ( w1029 , w1055 , w310 );
and ( w1030 , w1029 , w1064 );
and ( w1031 , w1030 , w13211 );
and ( w1032 , w1031 , w79 );
and ( w1033 , w1032 , w12612 );
nor ( w1034 , w1029 , w1033 );
nor ( w1035 , w1034 , w489 );
and ( w1036 , w1035 , w20 );
and ( w1037 , w1036 , w12080 );
and ( w1038 , w1037 , w8848 );
and ( w1039 , w1038 , w79 );
and ( w1040 , w1039 , w12612 );
nor ( w1041 , w1028 , w1040 );
nor ( w1042 , w713 , w632 );
not ( w1043 , w1042 );
and ( w1044 , w1043 , w310 );
and ( w1045 , w1044 , w377 );
and ( w1046 , w8848 , w649 );
and ( w1047 , w1046 , w255 );
and ( w1048 , w1047 , w20 );
not ( w1049 , w1048 );
and ( w1050 , w1049 , w626 );
not ( w1051 , w679 );
and ( w1052 , w1050 , w1051 );
not ( w1053 , w1052 );
and ( w1054 , w1053 , w312 );
not ( w1055 , w375 );
and ( w1056 , w798 , w1055 );
and ( w1057 , w1056 , w1231 );
and ( w1058 , w1057 , w8848 );
and ( w1059 , w1058 , w20 );
nor ( w1060 , w1059 , w634 );
not ( w1061 , w1060 );
and ( w1062 , w1061 , w377 );
nor ( w1063 , w1062 , w679 );
not ( w1064 , w309 );
and ( w1065 , w377 , w1064 );
and ( w1066 , w1065 , w13211 );
and ( w1067 , w1066 , w8848 );
and ( w1068 , w1067 , w20 );
and ( w1069 , w1068 , w79 );
and ( w1070 , w1069 , w12612 );
not ( w1071 , w1070 );
and ( w1072 , w1063 , w1071 );
and ( w1073 , w1072 , w12080 );
not ( w1074 , w1073 );
and ( w1075 , w1074 , w310 );
and ( w1076 , w1075 , w12080 );
and ( w1077 , w1076 , w310 );
and ( w1078 , w1077 , w79 );
and ( w1079 , w1078 , w12612 );
nor ( w1080 , w679 , w1079 );
nor ( w1081 , w19 , w383 );
and ( w1082 , w1081 , w20 );
not ( w1083 , w1082 );
and ( w1084 , w1083 , w626 );
nor ( w1085 , w309 , w383 );
and ( w1086 , w8848 , w1085 );
and ( w1087 , w1086 , w20 );
and ( w1088 , w1087 , w255 );
and ( w1089 , w1088 , w79 );
and ( w1090 , w1089 , w12612 );
not ( w1091 , w1090 );
and ( w1092 , w1084 , w1091 );
nor ( w1093 , w1092 , w648 );
and ( w1094 , w1093 , w255 );
and ( w1095 , w1094 , w11852 );
and ( w1096 , w1095 , w216 );
and ( w1097 , w1096 , w79 );
and ( w1098 , w1097 , w12612 );
not ( w1099 , w1098 );
and ( w1100 , w1080 , w1099 );
not ( w1101 , w1054 );
and ( w1102 , w1101 , w1100 );
nor ( w1103 , w1102 , w384 );
and ( w1104 , w1103 , w216 );
and ( w1105 , w1104 , w79 );
and ( w1106 , w1105 , w12612 );
nor ( w1107 , w1045 , w1106 );
not ( w1108 , w1107 );
and ( w1109 , w1108 , w312 );
not ( w1110 , w1109 );
and ( w1111 , w1110 , w1100 );
not ( w1112 , w1111 );
and ( w1113 , w1112 , w79 );
and ( w1114 , w1113 , w12612 );
not ( w1115 , w1114 );
and ( w1116 , w1041 , w1115 );
not ( w1117 , w1116 );
and ( w1118 , w1117 , w216 );
and ( w1119 , w1118 , w79 );
and ( w1120 , w1119 , w12612 );
nor ( w1121 , w1019 , w1120 );
not ( w1122 , w1121 );
and ( w1123 , w1122 , w79 );
nor ( w1124 , w1013 , w1123 );
and ( w1125 , w1124 , w111 );
and ( w1126 , w1125 , w125 );
nor ( w1127 , w1126 , w48 );
not ( w1128 , w1127 );
and ( w1129 , w1128 , w15 );
not ( w1130 , w1129 );
and ( w1131 , w1130 , w79 );
nor ( w1132 , w721 , w1131 );
not ( w1133 , w1123 );
and ( w1134 , w1132 , w1133 );
and ( w1135 , w1134 , w111 );
and ( w1136 , w1135 , w15 );
not ( w1137 , w1136 );
and ( w1138 , w1137 , w79 );
and ( w1139 , w1138 , w12612 );
not ( w1140 , w711 );
and ( w1141 , w1140 , w1139 );
not ( w1142 , w1141 );
and ( w1143 , w1142 , w15 );
not ( w1144 , w1143 );
and ( w1145 , w1144 , w79 );
and ( w1146 , w1145 , w12612 );
and ( w1147 , w701 , w1208 );
not ( w1148 , w1147 );
and ( w1149 , w1148 , w1139 );
nor ( w1150 , w1149 , w377 );
not ( w1151 , w1150 );
and ( w1152 , w1151 , g29 );
not ( w1153 , w1152 );
and ( w1154 , w1153 , g29 );
and ( w1155 , w1154 , w255 );
and ( w1156 , w553 , w8848 );
and ( w1157 , w1156 , w485 );
and ( w1158 , w1157 , w1452 );
nor ( w1159 , w1158 , w1146 );
and ( w1160 , w1159 , w12080 );
and ( w1161 , w12142 , w1160 );
and ( w1162 , w1161 , w125 );
nor ( w1163 , w1162 , w48 );
not ( w1164 , w1163 );
and ( w1165 , w1164 , w15 );
not ( w1166 , w1165 );
and ( w1167 , w1166 , w216 );
and ( w1168 , w1167 , w79 );
and ( w1169 , w1168 , w12612 );
not ( w1170 , w1155 );
and ( w1171 , w1170 , w1169 );
and ( w1172 , w1171 , w79 );
and ( w1173 , w1172 , w12612 );
nor ( w1174 , w485 , w1173 );
and ( w1175 , w1174 , w12921 );
and ( w1176 , w557 , w1452 );
nor ( w1177 , w1176 , w1139 );
and ( w1178 , w1177 , w8848 );
and ( w1179 , w1178 , w255 );
not ( w1180 , w1179 );
and ( w1181 , w1180 , w1169 );
and ( w1182 , w12142 , w1181 );
and ( w1183 , w1182 , w216 );
and ( w1184 , w1183 , w79 );
and ( w1185 , w1184 , w12612 );
and ( w1186 , w1185 , w1452 );
nor ( w1187 , w1186 , w1173 );
and ( w1188 , w1187 , w8848 );
and ( w1189 , w1188 , w12921 );
nor ( w1190 , w1189 , w489 );
and ( w1191 , w1190 , w1169 );
and ( w1192 , w1191 , w216 );
and ( w1193 , w1192 , w79 );
and ( w1194 , w1193 , w12612 );
and ( w1195 , w1194 , w485 );
nor ( w1196 , w1195 , w1173 );
and ( w1197 , w1196 , w8848 );
and ( w1198 , w1197 , w12921 );
nor ( w1199 , w1198 , w489 );
and ( w1200 , w1199 , w1169 );
and ( w1201 , w1200 , w79 );
and ( w1202 , w1201 , w12612 );
and ( w1203 , w1229 , w1202 );
and ( w1204 , w1203 , w1231 );
nor ( w1205 , w1204 , w19 );
nor ( w1206 , w679 , w632 );
and ( w1207 , w1206 , w105 );
not ( w1208 , w1146 );
and ( w1209 , w1207 , w1208 );
not ( w1210 , w1209 );
and ( w1211 , w1210 , w1139 );
not ( w1212 , w1211 );
and ( w1213 , w1212 , w486 );
and ( w1214 , w1213 , w19 );
and ( w1215 , w1214 , w12498 );
not ( w1216 , w1215 );
and ( w1217 , w1216 , g29 );
not ( w1218 , w1217 );
and ( w1219 , w1218 , g29 );
and ( w1220 , w1219 , w255 );
not ( w1221 , w1220 );
and ( w1222 , w1221 , w1169 );
and ( w1223 , w1222 , w79 );
and ( w1224 , w1223 , w12612 );
not ( w1225 , w1205 );
and ( w1226 , w1225 , w1224 );
and ( w1227 , w1226 , w79 );
and ( w1228 , w1227 , w12612 );
not ( w1229 , w1175 );
and ( w1230 , w1229 , w1228 );
not ( w1231 , w489 );
and ( w1232 , w1230 , w1231 );
not ( w1233 , w1139 );
and ( w1234 , w486 , w1233 );
nor ( w1235 , w1234 , w502 );
and ( w1236 , w1235 , w1224 );
and ( w1237 , w1236 , w216 );
and ( w1238 , w1237 , w12612 );
and ( w1239 , w1232 , w1238 );
nor ( w1240 , w1239 , w19 );
not ( w1241 , w1240 );
and ( w1242 , w1241 , w1224 );
and ( w1243 , w1242 , w79 );
and ( w1244 , w1243 , w12612 );
and ( w1245 , w700 , w1258 );
and ( w1246 , w1245 , w15 );
and ( w1247 , w1246 , w377 );
and ( w1248 , w1247 , w696 );
not ( w1249 , w1248 );
and ( w1250 , w1249 , w377 );
not ( w1251 , w1250 );
and ( w1252 , w1251 , w700 );
and ( w1253 , w1252 , w15 );
and ( w1254 , w686 , w1253 );
not ( w1255 , w1254 );
and ( w1256 , w19 , w1255 );
and ( w1257 , w1246 , w696 );
not ( w1258 , w1244 );
and ( w1259 , w1257 , w1258 );
and ( w1260 , w1259 , w15 );
not ( w1261 , w1256 );
and ( w1262 , w1261 , w1260 );
and ( w1263 , w1262 , w600 );
and ( w1264 , w1263 , w12921 );
nor ( w1265 , w1264 , w489 );
nor ( w1266 , w48 , w226 );
and ( w1267 , w1265 , w1278 );
nor ( w1268 , w1267 , w1244 );
and ( w1269 , w1268 , w15 );
not ( w1270 , w1269 );
and ( w1271 , w1270 , w216 );
and ( w1272 , w1271 , w79 );
and ( w1273 , w1272 , w12612 );
not ( w1274 , w674 );
and ( w1275 , w1274 , w1273 );
and ( w1276 , w1275 , w12919 );
and ( w1277 , w1276 , w48 );
not ( w1278 , w1266 );
and ( w1279 , w1277 , w1278 );
nor ( w1280 , w1279 , w1244 );
and ( w1281 , w1280 , w15 );
not ( w1282 , w1281 );
and ( w1283 , w1282 , w216 );
and ( w1284 , w1283 , w79 );
and ( w1285 , w1284 , w12612 );
not ( w1286 , w623 );
and ( w1287 , w1286 , w1285 );
and ( w1288 , w1287 , w216 );
and ( w1289 , w1288 , w79 );
not ( w1290 , w622 );
and ( w1291 , w1290 , w79 );
nor ( w1292 , w1289 , w1291 );
not ( w1293 , w1292 );
and ( w1294 , w1293 , w1285 );
not ( w1295 , w1294 );
and ( w1296 , w1295 , w15 );
not ( w1297 , w1296 );
and ( w1298 , w1297 , w216 );
and ( w1299 , w1298 , w79 );
nor ( w1300 , w1299 , w1291 );
and ( w1301 , w1300 , w19 );
nor ( w1302 , w1301 , w375 );
nor ( w1303 , w1302 , g12 );
and ( w1304 , w1303 , w111 );
and ( w1305 , w1304 , w11797 );
and ( w1306 , w1315 , w483 );
and ( w1307 , w1306 , w111 );
nor ( w1308 , w1307 , w105 );
not ( w1309 , w1308 );
and ( w1310 , w1309 , w125 );
nor ( w1311 , w1310 , w48 );
nor ( w1312 , w1311 , w19 );
not ( w1313 , w1299 );
and ( w1314 , w1313 , w483 );
not ( w1315 , w1291 );
and ( w1316 , w1314 , w1315 );
and ( w1317 , w1316 , w19 );
not ( w1318 , w1317 );
and ( w1319 , w1318 , w1285 );
not ( w1320 , w1319 );
and ( w1321 , w1320 , w15 );
not ( w1322 , w1321 );
and ( w1323 , w1322 , w216 );
and ( w1324 , w1323 , w79 );
not ( w1325 , w1312 );
and ( w1326 , w1325 , w1324 );
and ( w1327 , w1326 , w1285 );
not ( w1328 , w1327 );
and ( w1329 , w1328 , w15 );
not ( w1330 , w1329 );
and ( w1331 , w1330 , w216 );
and ( w1332 , w1331 , w79 );
and ( w1333 , w1332 , w12612 );
not ( w1334 , w1333 );
and ( w1335 , w1334 , w111 );
not ( w1336 , w661 );
and ( w1337 , w255 , w1336 );
not ( w1338 , w1337 );
and ( w1339 , w1338 , w108 );
and ( w1340 , w1339 , w12919 );
and ( w1341 , w1340 , w48 );
and ( w1342 , w536 , w485 );
and ( w1343 , w1342 , w12142 );
and ( w1344 , w1343 , w1452 );
and ( w1345 , w12142 , w1344 );
nor ( w1346 , w1345 , w20 );
nor ( w1347 , w1346 , w489 );
and ( w1348 , w1347 , w216 );
and ( w1349 , w1348 , w79 );
and ( w1350 , w1349 , w12612 );
and ( w1351 , w485 , w1350 );
nor ( w1352 , w1351 , w20 );
nor ( w1353 , w1352 , w489 );
and ( w1354 , w1353 , w79 );
and ( w1355 , w1354 , w12612 );
nor ( w1356 , w1341 , w1355 );
nor ( w1357 , w1356 , w105 );
not ( w1358 , w1357 );
and ( w1359 , w1358 , w600 );
nor ( w1360 , w621 , w1289 );
and ( w1361 , w1360 , w105 );
and ( w1362 , w1361 , w8640 );
and ( w1363 , w1362 , w522 );
and ( w1364 , w1363 , w105 );
and ( w1365 , w1364 , w8848 );
not ( w1366 , w1365 );
and ( w1367 , w1366 , w1285 );
not ( w1368 , w1367 );
and ( w1369 , w1368 , w15 );
not ( w1370 , w1369 );
and ( w1371 , w1370 , w216 );
and ( w1372 , w1371 , w79 );
and ( w1373 , w1372 , w12612 );
not ( w1374 , w1359 );
and ( w1375 , w1374 , w1373 );
and ( w1376 , w1375 , w1324 );
nor ( w1377 , w1376 , w20 );
nor ( w1378 , w1377 , w489 );
not ( w1379 , w1378 );
and ( w1380 , w1379 , w15 );
not ( w1381 , w1380 );
and ( w1382 , w1381 , w216 );
and ( w1383 , w1382 , w79 );
and ( w1384 , w1383 , w12612 );
not ( w1385 , w1384 );
and ( w1386 , w1335 , w1385 );
and ( w1387 , w1386 , w8848 );
not ( w1388 , w1387 );
and ( w1389 , w1388 , w1373 );
and ( w1390 , w1389 , w1324 );
nor ( w1391 , w1390 , w20 );
nor ( w1392 , w1391 , w489 );
not ( w1393 , w1392 );
and ( w1394 , w1393 , w15 );
not ( w1395 , w1394 );
and ( w1396 , w1395 , w216 );
and ( w1397 , w1396 , w79 );
and ( w1398 , w1397 , w12612 );
not ( w1399 , w1305 );
and ( w1400 , w1399 , w1398 );
and ( w1401 , w1400 , w1285 );
not ( w1402 , w1401 );
and ( w1403 , w1402 , w15 );
not ( w1404 , w1403 );
and ( w1405 , w1404 , w216 );
and ( w1406 , w1405 , w79 );
and ( w1407 , w1406 , w12612 );
not ( w1408 , w616 );
and ( w1409 , w1408 , w1407 );
and ( w1410 , w1409 , w1285 );
not ( w1411 , w1410 );
and ( w1412 , w1411 , w15 );
not ( w1413 , w1412 );
and ( w1414 , w1413 , w216 );
and ( w1415 , w1414 , w79 );
and ( w1416 , w1415 , w12612 );
not ( w1417 , w607 );
and ( w1418 , w1417 , w1416 );
nor ( w1419 , w1418 , w19 );
and ( w1420 , w1419 , w12921 );
nor ( w1421 , w1420 , w489 );
nor ( w1422 , w1421 , w312 );
not ( w1423 , w1422 );
and ( w1424 , w1423 , w1407 );
and ( w1425 , w1424 , w1285 );
not ( w1426 , w1425 );
and ( w1427 , w1426 , w15 );
not ( w1428 , w1427 );
and ( w1429 , w1428 , w216 );
and ( w1430 , w1429 , w79 );
and ( w1431 , w1430 , w12612 );
and ( w1432 , w602 , w1459 );
and ( w1433 , w1432 , w8848 );
and ( w1434 , w1433 , w12921 );
nor ( w1435 , w1434 , w489 );
not ( w1436 , w1435 );
and ( w1437 , w1436 , w15 );
not ( w1438 , w1437 );
and ( w1439 , w1438 , w216 );
and ( w1440 , w1439 , w79 );
and ( w1441 , w1440 , w12612 );
not ( w1442 , w1441 );
and ( w1443 , w586 , w1442 );
not ( w1444 , w1443 );
and ( w1445 , w1444 , w536 );
and ( w1446 , w12142 , w1445 );
not ( w1447 , w1446 );
and ( w1448 , w1447 , w483 );
and ( w1449 , w1448 , w12919 );
not ( w1450 , w1449 );
and ( w1451 , w1450 , w485 );
not ( w1452 , w486 );
and ( w1453 , w1451 , w1452 );
not ( w1454 , w1453 );
and ( w1455 , w1454 , w111 );
nor ( w1456 , w1455 , w105 );
not ( w1457 , w1456 );
and ( w1458 , w1457 , w600 );
not ( w1459 , w1431 );
and ( w1460 , w1458 , w1459 );
and ( w1461 , w1460 , w8848 );
and ( w1462 , w1461 , w12921 );
nor ( w1463 , w1462 , w489 );
and ( w1464 , w1463 , w1407 );
and ( w1465 , w1464 , w1285 );
not ( w1466 , w1465 );
and ( w1467 , w1466 , w15 );
not ( w1468 , w1467 );
and ( w1469 , w1468 , w216 );
and ( w1470 , w1469 , w79 );
and ( w1471 , w1470 , w12612 );
not ( w1472 , w488 );
and ( w1473 , w1472 , w1471 );
nor ( w1474 , w1473 , w20 );
nor ( w1475 , w1474 , w489 );
nor ( w1476 , w1475 , w312 );
not ( w1477 , w1476 );
and ( w1478 , w1477 , w1407 );
and ( w1479 , w1478 , w1285 );
not ( w1480 , w1479 );
and ( w1481 , w1480 , w15 );
not ( w1482 , w1481 );
and ( w1483 , w1482 , w216 );
and ( w1484 , w1483 , w79 );
and ( w1485 , w1484 , w12612 );
not ( w1486 , w406 );
and ( w1487 , w1486 , w1485 );
not ( w1488 , w1487 );
and ( w1489 , w1488 , w309 );
and ( w1490 , w1489 , w12037 );
not ( w1491 , w1490 );
and ( w1492 , w1491 , w1407 );
not ( w1493 , w1492 );
and ( w1494 , w1493 , w15 );
not ( w1495 , w1494 );
and ( w1496 , w1495 , w216 );
and ( w1497 , w1496 , w79 );
and ( w1498 , w1497 , w12612 );
nor ( w1499 , w398 , w1498 );
not ( w1500 , w1499 );
and ( w1501 , w1500 , w1485 );
and ( w1502 , w1501 , w1407 );
and ( w1503 , w1502 , w1285 );
and ( w1504 , w1503 , w216 );
and ( w1505 , w1504 , w79 );
and ( w1506 , w1505 , w12612 );
nor ( w1507 , w373 , w1506 );
and ( w1508 , w1507 , w17 );
nor ( w1509 , w1508 , w230 );
and ( w1510 , w1509 , w79 );
and ( w1511 , w1510 , w12612 );
not ( w1512 , w1511 );
and ( w1513 , w363 , w1512 );
nor ( w1514 , w18 , w1513 );
and ( w1515 , w12921 , w1514 );
not ( w1516 , w1515 );
and ( w1517 , w1516 , w111 );
and ( w1518 , w12921 , g12 );
not ( w1519 , w1518 );
and ( w1520 , w1519 , g13 );
not ( w1521 , w1520 );
and ( w1522 , w1521 , g13 );
nor ( w1523 , w1517 , w1522 );
nor ( w1524 , w1523 , w1506 );
and ( w1525 , w1524 , w17 );
and ( w1526 , w1525 , w15 );
nor ( w1527 , w1526 , w230 );
and ( w1528 , w1527 , w79 );
and ( w1529 , w1528 , w12612 );
nor ( w1530 , w307 , w1529 );
and ( w1531 , w1530 , w1607 );
and ( w1532 , w1531 , w17 );
nor ( w1533 , w1532 , w230 );
and ( w1534 , w1533 , w79 );
and ( w1535 , w1534 , w12612 );
not ( w1536 , w123 );
and ( w1537 , w1536 , w1535 );
and ( w1538 , w1537 , w12080 );
and ( w1539 , w1535 , w12080 );
nor ( w1540 , w383 , w380 );
and ( w1541 , w1540 , w255 );
not ( w1542 , w1541 );
and ( w1543 , w1542 , w17 );
not ( w1544 , w1539 );
and ( w1545 , w1544 , w1543 );
nor ( w1546 , w1545 , w309 );
not ( w1547 , w1546 );
and ( w1548 , w1547 , w308 );
nor ( w1549 , w1548 , w55 );
nor ( w1550 , w1549 , w304 );
nor ( w1551 , w20 , w1550 );
and ( w1552 , w8848 , w1551 );
nor ( w1553 , w1552 , w1529 );
and ( w1554 , w1553 , w1607 );
and ( w1555 , w1554 , w17 );
nor ( w1556 , w1555 , w230 );
and ( w1557 , w1556 , w79 );
and ( w1558 , w1557 , w12612 );
and ( w1559 , w1538 , w1558 );
not ( w1560 , w1559 );
and ( w1561 , w1560 , w1543 );
not ( w1562 , w1540 );
and ( w1563 , w255 , w1562 );
and ( w1564 , w1563 , w17 );
nor ( w1565 , w1564 , w255 );
nor ( w1566 , w1565 , w1540 );
and ( w1567 , w1566 , w17 );
nor ( w1568 , w1567 , w255 );
nor ( w1569 , w1568 , w1540 );
and ( w1570 , w1569 , w17 );
nor ( w1571 , w1561 , w1570 );
and ( w1572 , w1571 , w108 );
not ( w1573 , w103 );
and ( w1574 , w1572 , w1573 );
and ( w1575 , w1574 , w12919 );
nor ( w1576 , w1575 , w304 );
nor ( w1577 , w20 , w1576 );
and ( w1578 , w8848 , w1577 );
nor ( w1579 , w1578 , w1529 );
and ( w1580 , w1579 , w1607 );
and ( w1581 , w1580 , w17 );
nor ( w1582 , w1581 , w230 );
and ( w1583 , w1582 , w79 );
and ( w1584 , w1583 , w12612 );
and ( w1585 , w12919 , w1584 );
and ( w1586 , w1585 , w12921 );
nor ( w1587 , w1584 , w1511 );
and ( w1588 , w1587 , w12142 );
and ( w1589 , w1588 , w12921 );
nor ( w1590 , w1589 , w105 );
nor ( w1591 , w1590 , w485 );
nor ( w1592 , w1591 , w19 );
nor ( w1593 , w1592 , w1529 );
and ( w1594 , w1593 , w1607 );
and ( w1595 , w1594 , w17 );
nor ( w1596 , w1595 , w230 );
and ( w1597 , w1596 , w79 );
and ( w1598 , w1597 , w12612 );
and ( w1599 , w1586 , w1598 );
nor ( w1600 , w1599 , w1506 );
and ( w1601 , w1600 , w17 );
nor ( w1602 , w1601 , w230 );
and ( w1603 , w1602 , w216 );
and ( w1604 , w1603 , w79 );
and ( w1605 , w1604 , w12612 );
nor ( w1606 , w1605 , w1511 );
not ( w1607 , w1506 );
and ( w1608 , w1606 , w1607 );
and ( w1609 , w1608 , w17 );
nor ( w1610 , w1609 , w230 );
and ( w1611 , w1610 , w12612 );
and ( w1612 , w17 , w2393 );
and ( w1613 , w7 , w2501 );
nor ( w1614 , w1613 , w1611 );
nor ( w1615 , w1614 , w1612 );
nor ( w1616 , w1615 , g3 );
and ( w1617 , w1616 , w6138 );
nor ( w1618 , w1617 , w1612 );
and ( w1619 , w1618 , g5 );
and ( w1620 , w212 , w2501 );
nor ( w1621 , w1620 , w1615 );
not ( w1622 , w1619 );
and ( w1623 , w1622 , w1621 );
and ( w1624 , w1623 , w2396 );
and ( w1625 , w2396 , g36 );
nor ( w1626 , w73 , w1612 );
and ( w1627 , w1626 , g7 );
nor ( w1628 , w207 , g5 );
and ( w1629 , w1628 , w12934 );
and ( w1630 , w1629 , w2501 );
and ( w1631 , w1630 , w12934 );
and ( w1632 , w1626 , g5 );
nor ( w1633 , w1631 , w1632 );
not ( w1634 , w1627 );
and ( w1635 , w1634 , w1633 );
nor ( w1636 , w1625 , w1635 );
not ( w1637 , w1636 );
and ( w1638 , w1637 , g11 );
nor ( w1639 , w230 , w1612 );
nor ( w1640 , w1611 , w1615 );
and ( w1641 , g37 , w2501 );
and ( w1642 , w1641 , g19 );
nor ( w1643 , w1642 , w1615 );
and ( w1644 , w1640 , w1643 );
nor ( w1645 , w1644 , g19 );
not ( w1646 , w1645 );
and ( w1647 , w1640 , w1646 );
and ( w1648 , w1647 , w2396 );
and ( w1649 , w1648 , w1623 );
and ( w1650 , w1649 , w2396 );
and ( w1651 , w1650 , w1623 );
and ( w1652 , w1651 , w2396 );
and ( w1653 , w1652 , w1623 );
and ( w1654 , w1653 , w2396 );
and ( w1655 , w1654 , w1623 );
and ( w1656 , w1655 , w2396 );
and ( w1657 , w1656 , w1623 );
and ( w1658 , w1640 , w1657 );
and ( w1659 , w1658 , w2393 );
and ( w1660 , w1659 , w2396 );
and ( w1661 , w1658 , w1623 );
and ( w1662 , w1661 , w2396 );
and ( w1663 , w1662 , w1623 );
and ( w1664 , w1663 , w2396 );
and ( w1665 , w1664 , w1623 );
and ( w1666 , w1660 , w1665 );
and ( w1667 , g38 , w2501 );
and ( w1668 , w1667 , g25 );
nor ( w1669 , w1668 , w1615 );
and ( w1670 , w1666 , w1669 );
and ( w1671 , w2485 , g38 );
not ( w1672 , w1671 );
and ( w1673 , w1672 , g38 );
nor ( w1674 , w1673 , w1612 );
and ( w1675 , w1674 , g25 );
not ( w1676 , w1675 );
and ( w1677 , w1676 , g25 );
nor ( w1678 , w1670 , w1677 );
and ( w1679 , w2393 , g38 );
nor ( w1680 , w1679 , w1635 );
not ( w1681 , w1680 );
and ( w1682 , w1681 , g25 );
and ( w1683 , w1678 , w2126 );
and ( w1684 , w1624 , w1640 );
and ( w1685 , g39 , w2501 );
not ( w1686 , w1685 );
and ( w1687 , w1686 , g39 );
not ( w1688 , w1687 );
and ( w1689 , w1688 , g13 );
and ( w1690 , w1689 , w2485 );
not ( w1691 , w1690 );
and ( w1692 , w1691 , g13 );
nor ( w1693 , w1635 , g40 );
nor ( w1694 , w1693 , g40 );
nor ( w1695 , w1694 , w1612 );
and ( w1696 , w1695 , w9049 );
nor ( w1697 , w1696 , g17 );
not ( w1698 , w1697 );
and ( w1699 , w1698 , g15 );
and ( w1700 , w1699 , w2501 );
and ( w1701 , w1700 , g41 );
not ( w1702 , w1701 );
and ( w1703 , w1702 , g41 );
nor ( w1704 , w1703 , w1635 );
not ( w1705 , w1704 );
and ( w1706 , w1705 , g15 );
and ( w1707 , g40 , w2501 );
not ( w1708 , w1707 );
and ( w1709 , w1708 , g40 );
not ( w1710 , w1709 );
and ( w1711 , w1710 , g17 );
and ( w1712 , w1711 , w2485 );
not ( w1713 , w1712 );
and ( w1714 , w1713 , g17 );
nor ( w1715 , w1706 , w1714 );
and ( w1716 , w1715 , w2485 );
and ( w1717 , w1716 , w1639 );
and ( w1718 , w1717 , w2501 );
and ( w1719 , w1718 , w1639 );
and ( w1720 , w1719 , w2501 );
and ( w1721 , w1720 , w9195 );
nor ( w1722 , w1721 , g37 );
nor ( w1723 , w1722 , w1612 );
and ( w1724 , w1723 , g19 );
not ( w1725 , w1724 );
and ( w1726 , w1725 , g19 );
and ( w1727 , w1715 , w1639 );
and ( w1728 , w1727 , w2501 );
and ( w1729 , w1728 , w1639 );
and ( w1730 , w1729 , w2501 );
and ( w1731 , w1730 , w1639 );
and ( w1732 , w1731 , w2485 );
not ( w1733 , w1726 );
and ( w1734 , w1733 , w1732 );
and ( w1735 , w1734 , w2485 );
and ( w1736 , w1735 , w9354 );
and ( w1737 , w1736 , w1639 );
and ( w1738 , w1737 , w2501 );
nor ( w1739 , w1738 , g42 );
nor ( w1740 , w1739 , w1612 );
and ( w1741 , w1740 , w1639 );
and ( w1742 , w1741 , w2501 );
and ( w1743 , w1742 , g21 );
not ( w1744 , w1743 );
and ( w1745 , w1744 , g21 );
and ( w1746 , w1734 , w1639 );
and ( w1747 , w1746 , w2501 );
and ( w1748 , w1747 , w1639 );
and ( w1749 , w1748 , w2501 );
and ( w1750 , w1749 , g42 );
not ( w1751 , w1750 );
and ( w1752 , w1751 , g42 );
nor ( w1753 , w1752 , w1635 );
not ( w1754 , w1745 );
and ( w1755 , w1754 , w1753 );
and ( w1756 , w1755 , w1639 );
and ( w1757 , w1756 , w2501 );
and ( w1758 , g43 , w2501 );
not ( w1759 , w1758 );
and ( w1760 , w1759 , g43 );
not ( w1761 , w1760 );
and ( w1762 , w1761 , g23 );
and ( w1763 , w1762 , w2485 );
not ( w1764 , w1763 );
and ( w1765 , w1764 , g23 );
not ( w1766 , w1765 );
and ( w1767 , w1757 , w1766 );
and ( w1768 , w1767 , w1639 );
and ( w1769 , w1768 , w2501 );
and ( w1770 , w2485 , w1639 );
and ( w1771 , w1769 , w1770 );
not ( w1772 , w1667 );
and ( w1773 , w1772 , g38 );
not ( w1774 , w1773 );
and ( w1775 , w1774 , g25 );
and ( w1776 , w1775 , w2485 );
not ( w1777 , w1776 );
and ( w1778 , w1777 , g25 );
and ( w1779 , w1771 , w2423 );
and ( w1780 , w1779 , w1639 );
and ( w1781 , w1780 , w2501 );
and ( w1782 , g44 , w2501 );
not ( w1783 , w1782 );
and ( w1784 , w1783 , g44 );
not ( w1785 , w1784 );
and ( w1786 , w1785 , g27 );
and ( w1787 , w1786 , w2485 );
not ( w1788 , w1787 );
and ( w1789 , w1788 , g27 );
and ( w1790 , w1781 , w2426 );
and ( w1791 , w1790 , w1639 );
and ( w1792 , w1791 , w2501 );
and ( w1793 , w1792 , w1770 );
and ( w1794 , w1793 , w2501 );
and ( w1795 , w1794 , w2485 );
and ( w1796 , w1795 , w2501 );
and ( w1797 , w1796 , w1639 );
and ( w1798 , w2488 , w1797 );
and ( w1799 , w1798 , w1639 );
and ( w1800 , w1799 , w2501 );
and ( w1801 , w1800 , w1639 );
and ( w1802 , w1801 , w2485 );
and ( w1803 , w1802 , w13474 );
and ( w1804 , w1803 , w13477 );
nor ( w1805 , w1804 , w1611 );
and ( w1806 , w1639 , w11795 );
and ( w1807 , w1806 , w11797 );
nor ( w1808 , w1807 , w1611 );
and ( w1809 , w1805 , w1808 );
not ( w1810 , w1809 );
and ( w1811 , w1810 , w1639 );
and ( w1812 , w1811 , w2485 );
and ( w1813 , w1812 , w1639 );
and ( w1814 , w1813 , w2485 );
and ( w1815 , w1814 , w13331 );
and ( w1816 , w1815 , w13333 );
nor ( w1817 , w1816 , w1615 );
and ( w1818 , w2393 , g36 );
nor ( w1819 , w1818 , w1635 );
not ( w1820 , w1819 );
and ( w1821 , w1820 , g11 );
nor ( w1822 , w1817 , w1821 );
nor ( w1823 , w1822 , w1611 );
and ( w1824 , w1823 , w2396 );
and ( w1825 , w1824 , w1623 );
and ( w1826 , w2393 , w1623 );
and ( w1827 , w1825 , w1826 );
and ( w1828 , w1684 , w1827 );
and ( w1829 , w1798 , w2485 );
and ( w1830 , w1829 , w1639 );
and ( w1831 , w1830 , w2501 );
and ( w1832 , w1831 , g45 );
and ( w1833 , w1832 , g29 );
nor ( w1834 , w1833 , w1611 );
nor ( w1835 , w1834 , g11 );
not ( w1836 , w1835 );
and ( w1837 , w1836 , w1808 );
not ( w1838 , w1837 );
and ( w1839 , w1838 , w1639 );
and ( w1840 , w1839 , w2522 );
and ( w1841 , w1840 , w1639 );
and ( w1842 , w1841 , w2485 );
and ( w1843 , w1842 , w13474 );
nor ( w1844 , w1843 , w1611 );
and ( w1845 , w1844 , w1808 );
not ( w1846 , w1845 );
and ( w1847 , w1846 , w1639 );
and ( w1848 , w2485 , g45 );
and ( w1849 , w1848 , g29 );
nor ( w1850 , w1849 , w1611 );
and ( w1851 , w1850 , w11795 );
and ( w1852 , w1851 , w11797 );
and ( w1853 , g39 , g13 );
and ( w1854 , w1852 , w13545 );
nor ( w1855 , w1854 , w1612 );
nor ( w1856 , w1855 , w1611 );
not ( w1857 , w1856 );
and ( w1858 , w1857 , w1639 );
and ( w1859 , w1858 , w2501 );
and ( w1860 , w1859 , w1639 );
and ( w1861 , w1860 , w2485 );
and ( w1862 , w1861 , w1639 );
and ( w1863 , w1847 , w1862 );
not ( w1864 , w1863 );
and ( w1865 , w1864 , w1640 );
not ( w1866 , w1822 );
and ( w1867 , w1865 , w1866 );
nor ( w1868 , w1867 , w1821 );
and ( w1869 , w1828 , w2504 );
not ( w1870 , w1683 );
and ( w1871 , w1870 , w1869 );
and ( w1872 , w1871 , w1826 );
and ( w1873 , w1872 , w1624 );
nor ( w1874 , g46 , w1612 );
and ( w1875 , w1874 , w13590 );
nor ( w1876 , w1875 , w1615 );
and ( w1877 , w1640 , w1876 );
nor ( w1878 , g46 , g9 );
nor ( w1879 , w1878 , w17 );
not ( w1880 , w1877 );
and ( w1881 , w1880 , w1879 );
nor ( w1882 , w1881 , w1611 );
and ( w1883 , w1882 , w1640 );
and ( w1884 , w1883 , w2393 );
and ( w1885 , w1884 , w1640 );
and ( w1886 , w1885 , w2393 );
and ( w1887 , w1886 , w1638 );
and ( w1888 , w1887 , w1821 );
and ( w1889 , w1640 , w1876 );
not ( w1890 , w1889 );
and ( w1891 , w1890 , w1879 );
nor ( w1892 , w1891 , w1611 );
and ( w1893 , w1892 , w1640 );
and ( w1894 , w1893 , w2393 );
and ( w1895 , w1894 , w1638 );
and ( w1896 , w1895 , w1821 );
and ( w1897 , w1624 , w1876 );
and ( w1898 , w1897 , w1640 );
not ( w1899 , w1898 );
and ( w1900 , w1899 , w1879 );
nor ( w1901 , w1900 , w1611 );
and ( w1902 , w1901 , w1826 );
nor ( w1903 , w1635 , g44 );
and ( w1904 , w1903 , w13050 );
not ( w1905 , w1904 );
and ( w1906 , w1905 , w1623 );
and ( w1907 , w1902 , w1906 );
nor ( w1908 , w1635 , g46 );
and ( w1909 , w1908 , w13590 );
not ( w1910 , w1909 );
and ( w1911 , w1910 , w1623 );
and ( w1912 , w1907 , w1911 );
and ( w1913 , w1912 , w2396 );
and ( w1914 , w1913 , w1623 );
nor ( w1915 , w1896 , w1914 );
and ( w1916 , w1888 , w1928 );
nor ( w1917 , w1916 , w1914 );
nor ( w1918 , w1917 , w1615 );
and ( w1919 , w1918 , w1623 );
and ( w1920 , w1873 , w1919 );
and ( w1921 , w1827 , w1682 );
nor ( w1922 , w1921 , w1677 );
not ( w1923 , w1669 );
and ( w1924 , w1922 , w1923 );
not ( w1925 , w1924 );
and ( w1926 , w1925 , w1826 );
and ( w1927 , w1926 , w1624 );
not ( w1928 , w1915 );
and ( w1929 , w1927 , w1928 );
and ( w1930 , w1929 , w1640 );
and ( w1931 , w1930 , w2393 );
nor ( w1932 , w1931 , w1612 );
and ( w1933 , w1932 , w2485 );
and ( w1934 , g46 , g9 );
not ( w1935 , w17 );
and ( w1936 , w1934 , w1935 );
nor ( w1937 , w1933 , w1936 );
and ( w1938 , w1937 , w2393 );
and ( w1939 , w1938 , w1624 );
and ( w1940 , w1623 , g46 );
nor ( w1941 , w1940 , w1612 );
not ( w1942 , w1941 );
and ( w1943 , w1942 , g9 );
nor ( w1944 , w1939 , w1943 );
not ( w1945 , w1944 );
and ( w1946 , w1945 , w1827 );
and ( w1947 , w1640 , w1876 );
not ( w1948 , w1947 );
and ( w1949 , w1948 , w1879 );
nor ( w1950 , w1949 , w1611 );
and ( w1951 , w2396 , g39 );
nor ( w1952 , w1951 , w1635 );
not ( w1953 , w1952 );
and ( w1954 , w1953 , g13 );
and ( w1955 , w1640 , w1638 );
and ( w1956 , w1623 , g41 );
nor ( w1957 , w1956 , w1635 );
not ( w1958 , w1957 );
and ( w1959 , w1958 , g15 );
and ( w1960 , w1623 , g37 );
nor ( w1961 , w1960 , w1635 );
not ( w1962 , w1961 );
and ( w1963 , w1962 , g19 );
nor ( w1964 , w1959 , w1963 );
and ( w1965 , w1959 , g37 );
nor ( w1966 , w1965 , w1635 );
not ( w1967 , w1641 );
and ( w1968 , w1967 , g37 );
not ( w1969 , w1968 );
and ( w1970 , w1969 , g19 );
and ( w1971 , w1970 , w2485 );
not ( w1972 , w1971 );
and ( w1973 , w1972 , g19 );
not ( w1974 , w1973 );
and ( w1975 , w1966 , w1974 );
and ( w1976 , w1975 , w9197 );
nor ( w1977 , w1964 , w1976 );
and ( w1978 , w2396 , g40 );
nor ( w1979 , w1978 , w1635 );
not ( w1980 , w1979 );
and ( w1981 , w1980 , g17 );
nor ( w1982 , w1977 , w1981 );
not ( w1983 , w1982 );
and ( w1984 , w1983 , w1624 );
and ( w1985 , w1693 , w9049 );
nor ( w1986 , w1985 , w1615 );
and ( w1987 , w1984 , w1986 );
nor ( w1988 , w1987 , w1963 );
nor ( w1989 , w1988 , w1615 );
and ( w1990 , w1989 , w1623 );
and ( w1991 , w1990 , w2396 );
and ( w1992 , w1991 , w1623 );
nor ( w1993 , w1635 , g37 );
and ( w1994 , w1993 , w9197 );
nor ( w1995 , w1994 , w1615 );
and ( w1996 , w1992 , w1995 );
nor ( w1997 , w1635 , g42 );
and ( w1998 , w1997 , w9356 );
not ( w1999 , w1998 );
and ( w2000 , w1999 , w1623 );
and ( w2001 , w1996 , w2000 );
and ( w2002 , w1623 , g42 );
nor ( w2003 , w2002 , w1635 );
not ( w2004 , w2003 );
and ( w2005 , w2004 , g21 );
nor ( w2006 , w2001 , w2005 );
nor ( w2007 , w2006 , w1615 );
and ( w2008 , w2007 , w1623 );
nor ( w2009 , w1635 , g43 );
and ( w2010 , w2009 , w13321 );
not ( w2011 , w2010 );
and ( w2012 , w2011 , w1623 );
and ( w2013 , w2008 , w2012 );
and ( w2014 , w1623 , g38 );
nor ( w2015 , w2014 , w1635 );
not ( w2016 , w2015 );
and ( w2017 , w2016 , g25 );
nor ( w2018 , w2013 , w2017 );
and ( w2019 , w1623 , g43 );
nor ( w2020 , w2019 , w1635 );
not ( w2021 , w2020 );
and ( w2022 , w2021 , g23 );
not ( w2023 , w2022 );
and ( w2024 , w2018 , w2023 );
nor ( w2025 , w2024 , w1615 );
and ( w2026 , w2025 , w1623 );
nor ( w2027 , w1635 , g38 );
and ( w2028 , w2027 , w12964 );
not ( w2029 , w2028 );
and ( w2030 , w2029 , w1623 );
and ( w2031 , w2026 , w2030 );
and ( w2032 , w2393 , g44 );
nor ( w2033 , w2032 , w1635 );
not ( w2034 , w2033 );
and ( w2035 , w2034 , g27 );
nor ( w2036 , w2031 , w2035 );
not ( w2037 , w2036 );
and ( w2038 , w2037 , w1640 );
and ( w2039 , w2038 , w1876 );
and ( w2040 , w2039 , w1624 );
and ( w2041 , w2040 , w1640 );
not ( w2042 , w2041 );
and ( w2043 , w2042 , w1879 );
nor ( w2044 , w2043 , w1611 );
and ( w2045 , w2044 , w1826 );
and ( w2046 , w2045 , w1906 );
and ( w2047 , w2046 , w1911 );
nor ( w2048 , w2047 , w1612 );
and ( w2049 , w2048 , w2485 );
and ( w2050 , w2049 , w2261 );
nor ( w2051 , w2050 , w1615 );
and ( w2052 , w2051 , w1623 );
and ( w2053 , w1684 , w1869 );
and ( w2054 , w2053 , w2504 );
and ( w2055 , w2054 , w1826 );
and ( w2056 , w2485 , g44 );
and ( w2057 , w2056 , g27 );
not ( w2058 , w2057 );
and ( w2059 , w2058 , w1623 );
nor ( w2060 , w2035 , w2059 );
not ( w2061 , w2060 );
and ( w2062 , w2061 , w1826 );
and ( w2063 , w2055 , w2062 );
and ( w2064 , w2063 , w1826 );
and ( w2065 , w2052 , w2064 );
and ( w2066 , w2065 , w1624 );
and ( w2067 , w2485 , g39 );
and ( w2068 , w2067 , g13 );
not ( w2069 , w2068 );
and ( w2070 , w2069 , w1623 );
and ( w2071 , w2066 , w2070 );
and ( w2072 , w2071 , w1624 );
nor ( w2073 , w1635 , g36 );
and ( w2074 , w2073 , w13477 );
not ( w2075 , w2074 );
and ( w2076 , w2075 , w1623 );
and ( w2077 , w2072 , w2076 );
nor ( w2078 , w1955 , w2077 );
nor ( w2079 , w2078 , w1611 );
nor ( w2080 , w2079 , w1635 );
and ( w2081 , w2080 , w13331 );
and ( w2082 , w2081 , w13333 );
nor ( w2083 , w2082 , w1615 );
nor ( w2084 , w1683 , w1868 );
and ( w2085 , w2084 , w1640 );
and ( w2086 , w2085 , w2396 );
and ( w2087 , w2086 , w1623 );
and ( w2088 , w1624 , w1986 );
nor ( w2089 , w2088 , w1963 );
not ( w2090 , w2089 );
and ( w2091 , w2090 , w1995 );
and ( w2092 , w2091 , w2000 );
and ( w2093 , g42 , w2501 );
and ( w2094 , w2093 , g21 );
nor ( w2095 , w2094 , w1615 );
and ( w2096 , w2092 , w2095 );
and ( w2097 , w2096 , w2001 );
not ( w2098 , w2097 );
and ( w2099 , w2098 , w1639 );
and ( w2100 , w2099 , w2501 );
and ( w2101 , w2100 , w1770 );
and ( w2102 , w2101 , w2311 );
not ( w2103 , w2102 );
and ( w2104 , w2103 , w1624 );
nor ( w2105 , w2104 , w2022 );
not ( w2106 , w2105 );
and ( w2107 , w2106 , w2012 );
and ( w2108 , w2107 , w2030 );
nor ( w2109 , w2108 , w2035 );
not ( w2110 , w2109 );
and ( w2111 , w2110 , w1640 );
and ( w2112 , w2111 , w1624 );
nor ( w2113 , w2112 , w2017 );
nor ( w2114 , w2113 , w1615 );
and ( w2115 , w2114 , w1623 );
and ( w2116 , w2115 , w2064 );
and ( w2117 , w2116 , w1624 );
and ( w2118 , w2087 , w2117 );
and ( w2119 , w2118 , w1640 );
and ( w2120 , w2119 , w1826 );
and ( w2121 , w2120 , w1906 );
and ( w2122 , w2121 , w1911 );
and ( w2123 , w1640 , w1666 );
and ( w2124 , w2123 , w1669 );
nor ( w2125 , w2124 , w1677 );
not ( w2126 , w1682 );
and ( w2127 , w2125 , w2126 );
not ( w2128 , w2127 );
and ( w2129 , w2128 , w1826 );
and ( w2130 , w2129 , w1624 );
and ( w2131 , w2130 , w2396 );
and ( w2132 , w2131 , w1623 );
and ( w2133 , w1624 , w2095 );
not ( w2134 , w2133 );
and ( w2135 , w2134 , w1639 );
and ( w2136 , w2135 , w2501 );
and ( w2137 , w2136 , w1770 );
and ( w2138 , w2137 , w2311 );
not ( w2139 , w2138 );
and ( w2140 , w2139 , w1624 );
and ( w2141 , w2140 , w1638 );
and ( w2142 , w1623 , g40 );
nor ( w2143 , w2142 , w1635 );
not ( w2144 , w2143 );
and ( w2145 , w2144 , g17 );
and ( w2146 , w1624 , w2145 );
nor ( w2147 , w2146 , w1977 );
not ( w2148 , w2147 );
and ( w2149 , w2148 , w1624 );
and ( w2150 , w2149 , w1986 );
nor ( w2151 , w2150 , w1963 );
not ( w2152 , w2151 );
and ( w2153 , w2152 , w2000 );
and ( w2154 , w2153 , w1995 );
nor ( w2155 , w2154 , w2005 );
not ( w2156 , w2155 );
and ( w2157 , w2156 , w2012 );
nor ( w2158 , w2157 , w2022 );
not ( w2159 , w2158 );
and ( w2160 , w2159 , w2030 );
nor ( w2161 , w2160 , w1682 );
not ( w2162 , w2035 );
and ( w2163 , w2161 , w2162 );
not ( w2164 , w2163 );
and ( w2165 , w2164 , w1640 );
and ( w2166 , w2165 , w1624 );
and ( w2167 , w2166 , w1826 );
and ( w2168 , w2167 , w1911 );
and ( w2169 , w2168 , w1826 );
and ( w2170 , w2169 , w1906 );
and ( w2171 , w2485 , g36 );
and ( w2172 , w2171 , g11 );
not ( w2173 , w2172 );
and ( w2174 , w2173 , w1623 );
and ( w2175 , w2174 , w13331 );
nor ( w2176 , w2175 , w1635 );
and ( w2177 , w2176 , g29 );
not ( w2178 , w2174 );
and ( w2179 , w2178 , g45 );
not ( w2180 , w2179 );
and ( w2181 , w2180 , w1623 );
not ( w2182 , w2177 );
and ( w2183 , w2182 , w2181 );
nor ( w2184 , w2170 , w2183 );
nor ( w2185 , w2184 , w1868 );
and ( w2186 , w2185 , w2393 );
and ( w2187 , w2186 , g45 );
nor ( w2188 , w2187 , w1635 );
not ( w2189 , w2183 );
and ( w2190 , w2188 , w2189 );
not ( w2191 , w2190 );
and ( w2192 , w2191 , w2181 );
and ( w2193 , w2192 , w1640 );
and ( w2194 , w2193 , w1624 );
nor ( w2195 , w2141 , w2194 );
not ( w2196 , w2195 );
and ( w2197 , w2196 , w1624 );
and ( w2198 , w2197 , w2064 );
and ( w2199 , w2198 , w2070 );
and ( w2200 , w2132 , w2199 );
and ( w2201 , w2200 , w1826 );
and ( w2202 , w2201 , w1624 );
and ( w2203 , w2202 , w2504 );
and ( w2204 , w2203 , w1826 );
and ( w2205 , w2204 , w1638 );
and ( w2206 , w2205 , w1821 );
nor ( w2207 , w2206 , w1954 );
not ( w2208 , w2207 );
and ( w2209 , w2208 , w1640 );
nor ( w2210 , w2209 , w1612 );
and ( w2211 , w2210 , w2485 );
not ( w2212 , w2211 );
and ( w2213 , w2212 , w1624 );
nor ( w2214 , w2213 , w1943 );
not ( w2215 , w2214 );
and ( w2216 , w2215 , w1826 );
and ( w2217 , w2216 , w2504 );
and ( w2218 , w2217 , w1826 );
nor ( w2219 , w2122 , w2218 );
not ( w2220 , w2219 );
and ( w2221 , w2220 , w2070 );
nor ( w2222 , w2221 , w1954 );
not ( w2223 , w2222 );
and ( w2224 , w2223 , w1640 );
nor ( w2225 , w2224 , w1612 );
and ( w2226 , w2225 , w2485 );
and ( w2227 , w2226 , w2261 );
not ( w2228 , w2227 );
and ( w2229 , w2228 , w1826 );
and ( w2230 , w2229 , w2504 );
and ( w2231 , w2230 , w1624 );
and ( w2232 , w1623 , g45 );
nor ( w2233 , w2232 , w1635 );
not ( w2234 , w2233 );
and ( w2235 , w2234 , g29 );
nor ( w2236 , w2235 , w2077 );
not ( w2237 , w2236 );
and ( w2238 , w2237 , w1914 );
and ( w2239 , w2396 , g46 );
nor ( w2240 , w2239 , w1635 );
not ( w2241 , w2240 );
and ( w2242 , w2241 , g9 );
nor ( w2243 , w2238 , w2242 );
nor ( w2244 , g45 , w1635 );
nor ( w2245 , w2244 , w1615 );
nor ( w2246 , w2245 , w2183 );
not ( w2247 , w2246 );
and ( w2248 , w2247 , w2181 );
not ( w2249 , w2243 );
and ( w2250 , w2249 , w2248 );
and ( w2251 , w2198 , w2396 );
and ( w2252 , w2251 , w1623 );
and ( w2253 , w2252 , w2396 );
and ( w2254 , w2253 , w1623 );
and ( w2255 , w2254 , w1640 );
and ( w2256 , w2255 , w1826 );
and ( w2257 , w2256 , w1906 );
nor ( w2258 , w2257 , w2183 );
and ( w2259 , w2258 , w2501 );
and ( w2260 , w2259 , w2485 );
not ( w2261 , w1943 );
and ( w2262 , w2260 , w2261 );
not ( w2263 , w2262 );
and ( w2264 , w2263 , w1826 );
and ( w2265 , w2264 , w2504 );
and ( w2266 , w2265 , w1876 );
and ( w2267 , w2266 , w2393 );
not ( w2268 , w2267 );
and ( w2269 , w2268 , w1879 );
nor ( w2270 , w2269 , w1611 );
and ( w2271 , w2270 , w1826 );
and ( w2272 , w2271 , w1911 );
nor ( w2273 , w2272 , w2183 );
nor ( w2274 , w2273 , w1615 );
and ( w2275 , w2274 , w1624 );
and ( w2276 , w2275 , w2070 );
nor ( w2277 , w2276 , w1954 );
not ( w2278 , w2277 );
and ( w2279 , w2278 , w1624 );
and ( w2280 , w2250 , w2279 );
nor ( w2281 , w2280 , w1954 );
and ( w2282 , w2281 , w2491 );
not ( w2283 , w2282 );
and ( w2284 , w2283 , w1640 );
and ( w2285 , w2284 , w1624 );
and ( w2286 , w2285 , w2076 );
and ( w2287 , w2231 , w2286 );
and ( w2288 , w2287 , w1640 );
and ( w2289 , w2288 , w1826 );
and ( w2290 , w2289 , w2076 );
and ( w2291 , w2083 , w2290 );
nor ( w2292 , w1954 , w2291 );
not ( w2293 , w2292 );
and ( w2294 , w1950 , w2293 );
and ( w2295 , w2294 , w2393 );
not ( w2296 , w1936 );
and ( w2297 , w2295 , w2296 );
and ( w2298 , w2297 , w2393 );
and ( w2299 , w2298 , w1821 );
nor ( w2300 , w2299 , w1943 );
not ( w2301 , w2077 );
and ( w2302 , w2300 , w2301 );
not ( w2303 , w2302 );
and ( w2304 , w2303 , w1640 );
and ( w2305 , w1624 , w2064 );
and ( w2306 , w1624 , w2095 );
not ( w2307 , w2306 );
and ( w2308 , w2307 , w1639 );
and ( w2309 , w2308 , w2501 );
and ( w2310 , w2309 , w1770 );
not ( w2311 , w2005 );
and ( w2312 , w2310 , w2311 );
not ( w2313 , w2312 );
and ( w2314 , w2313 , w1624 );
and ( w2315 , w2305 , w2314 );
and ( w2316 , w2304 , w2315 );
and ( w2317 , w2316 , w2064 );
and ( w2318 , w2317 , w2314 );
and ( w2319 , w2318 , w1624 );
and ( w2320 , w2319 , w2393 );
nor ( w2321 , w2320 , w1692 );
nor ( w2322 , w2321 , w1853 );
nor ( w2323 , w2322 , w1612 );
nor ( w2324 , w2323 , w1611 );
and ( w2325 , w1623 , g39 );
nor ( w2326 , w2325 , w1612 );
not ( w2327 , w2326 );
and ( w2328 , w2327 , g13 );
nor ( w2329 , w2324 , w2328 );
and ( w2330 , w1826 , g39 );
nor ( w2331 , w2330 , w1635 );
not ( w2332 , w2331 );
and ( w2333 , w2332 , g13 );
and ( w2334 , w1827 , w2333 );
and ( w2335 , w2334 , w1640 );
and ( w2336 , w2335 , w1954 );
nor ( w2337 , w2336 , w2070 );
not ( w2338 , w2337 );
and ( w2339 , w2338 , w1826 );
not ( w2340 , w2329 );
and ( w2341 , w2340 , w2339 );
nor ( w2342 , w2341 , w1635 );
nor ( w2343 , w2342 , w1611 );
nor ( w2344 , w2343 , g45 );
and ( w2345 , w2344 , w13333 );
not ( w2346 , w2345 );
and ( w2347 , w2346 , w1826 );
and ( w2348 , w2347 , w2396 );
and ( w2349 , w2348 , w1624 );
and ( w2350 , w2349 , w2290 );
and ( w2351 , w2350 , w1624 );
and ( w2352 , w2351 , w2076 );
and ( w2353 , w1946 , w2352 );
and ( w2354 , w2353 , w2393 );
nor ( w2355 , w2354 , w1692 );
nor ( w2356 , w2355 , w1853 );
nor ( w2357 , w2356 , w1612 );
nor ( w2358 , w2357 , w1611 );
and ( w2359 , w2358 , w1624 );
nor ( w2360 , w2359 , w2328 );
not ( w2361 , w2360 );
and ( w2362 , w2361 , w2339 );
and ( w2363 , w2362 , w2393 );
and ( w2364 , w2363 , w1826 );
and ( w2365 , w2364 , w2396 );
and ( w2366 , w2365 , w1624 );
and ( w2367 , w2366 , w2290 );
and ( w2368 , w2367 , w1624 );
and ( w2369 , w2368 , w2076 );
and ( w2370 , w1920 , w2369 );
and ( w2371 , w2370 , w2393 );
nor ( w2372 , w2371 , w1612 );
and ( w2373 , w2372 , w2485 );
nor ( w2374 , w2373 , w1936 );
and ( w2375 , w2374 , w2393 );
and ( w2376 , w2375 , w1624 );
nor ( w2377 , w2376 , w1943 );
not ( w2378 , w2377 );
and ( w2379 , w2378 , w1827 );
and ( w2380 , w2379 , w1640 );
and ( w2381 , w2380 , w2396 );
and ( w2382 , w2381 , w1623 );
and ( w2383 , w2382 , w2352 );
and ( w2384 , w2383 , w2393 );
nor ( w2385 , w2384 , w1692 );
nor ( w2386 , w2385 , w1853 );
nor ( w2387 , w2386 , w1612 );
nor ( w2388 , w2387 , w1611 );
and ( w2389 , w2388 , w1624 );
nor ( w2390 , w2389 , w2328 );
not ( w2391 , w2390 );
and ( w2392 , w2391 , w2339 );
not ( w2393 , w1611 );
and ( w2394 , w2392 , w2393 );
and ( w2395 , w2394 , w1826 );
not ( w2396 , w1615 );
and ( w2397 , w2395 , w2396 );
and ( w2398 , w2397 , w1624 );
and ( w2399 , w2398 , w2290 );
and ( w2400 , w2399 , w1826 );
and ( w2401 , w2400 , w1624 );
and ( w2402 , w2401 , w2076 );
nor ( w2403 , g39 , w1612 );
and ( w2404 , w2403 , w11797 );
not ( w2405 , w2404 );
and ( w2406 , w2405 , w1623 );
and ( w2407 , w2402 , w2406 );
and ( w2408 , w2407 , w1808 );
nor ( w2409 , w2403 , g39 );
nor ( w2410 , w2409 , g13 );
and ( w2411 , w2410 , w2485 );
nor ( w2412 , w2411 , g13 );
nor ( w2413 , w2408 , w2412 );
and ( w2414 , w1770 , w1797 );
and ( w2415 , w2414 , w2501 );
and ( w2416 , w2415 , w2485 );
and ( w2417 , w2416 , w2501 );
and ( w2418 , w2417 , w1639 );
and ( w2419 , w1770 , w2418 );
and ( w2420 , w2419 , w2488 );
and ( w2421 , w2420 , w1639 );
and ( w2422 , w2421 , w2501 );
not ( w2423 , w1778 );
and ( w2424 , w2423 , w1639 );
and ( w2425 , w2424 , w2501 );
not ( w2426 , w1789 );
and ( w2427 , w2425 , w2426 );
and ( w2428 , w2427 , w1639 );
and ( w2429 , w2428 , w2501 );
and ( w2430 , w1770 , w2429 );
and ( w2431 , w2422 , w2430 );
and ( w2432 , w2431 , w1770 );
and ( w2433 , w2430 , w2488 );
and ( w2434 , w2433 , w1639 );
and ( w2435 , w2434 , w2501 );
and ( w2436 , w2435 , w2485 );
and ( w2437 , w2436 , w2501 );
and ( w2438 , w2437 , w1639 );
and ( w2439 , g36 , w2501 );
not ( w2440 , w2439 );
and ( w2441 , w2440 , g36 );
not ( w2442 , w2441 );
and ( w2443 , w2442 , g11 );
and ( w2444 , w2443 , w2485 );
not ( w2445 , w2444 );
and ( w2446 , w2445 , g11 );
and ( w2447 , w2438 , w2466 );
and ( w2448 , w2447 , w2488 );
and ( w2449 , w2448 , w1639 );
and ( w2450 , w2449 , w2501 );
and ( w2451 , w2450 , w2485 );
and ( w2452 , w2451 , w1639 );
and ( w2453 , w2452 , w2501 );
and ( w2454 , w2453 , w1639 );
and ( w2455 , w2454 , w2475 );
and ( w2456 , w2455 , w1639 );
and ( w2457 , w2456 , w2501 );
and ( w2458 , w2457 , w2466 );
and ( w2459 , w2458 , w2488 );
and ( w2460 , w2459 , w1639 );
and ( w2461 , w2460 , w2501 );
and ( w2462 , w2461 , w2485 );
and ( w2463 , w2462 , w1639 );
and ( w2464 , w2463 , w2501 );
and ( w2465 , w2464 , w1639 );
not ( w2466 , w2446 );
and ( w2467 , w2465 , w2466 );
and ( w2468 , w2467 , w2488 );
and ( w2469 , w2468 , w1639 );
and ( w2470 , w2469 , w2501 );
and ( w2471 , w2470 , w2485 );
and ( w2472 , w2471 , w1639 );
and ( w2473 , w2472 , w2501 );
and ( w2474 , w2473 , w1639 );
not ( w2475 , w2412 );
and ( w2476 , w2474 , w2475 );
and ( w2477 , w2476 , w1639 );
and ( w2478 , w2477 , w2501 );
and ( w2479 , w2432 , w2478 );
and ( w2480 , w1770 , w2479 );
and ( w2481 , w2413 , w2480 );
and ( w2482 , w2481 , w1639 );
and ( w2483 , w2482 , w2501 );
and ( w2484 , w1639 , w2483 );
not ( w2485 , w1635 );
and ( w2486 , w2484 , w2485 );
and ( w2487 , w2484 , w2501 );
not ( w2488 , w1692 );
and ( w2489 , w2488 , w2487 );
and ( w2490 , w2486 , w2489 );
not ( w2491 , w1638 );
and ( w2492 , w2491 , w2490 );
and ( w2493 , w1624 , w2183 );
not ( w2494 , w2493 );
and ( w2495 , w2494 , w2490 );
and ( w2496 , w2495 , w2489 );
and ( w2497 , w2496 , w2486 );
and ( w2498 , w2497 , w2490 );
and ( w2499 , w2498 , w2522 );
and ( w2500 , w1853 , w2487 );
not ( w2501 , w1612 );
and ( w2502 , w2500 , w2501 );
nor ( w2503 , w2502 , w1611 );
not ( w2504 , w1868 );
and ( w2505 , w2504 , w2503 );
and ( w2506 , g39 , w2484 );
nor ( w2507 , w2506 , w1611 );
and ( w2508 , g13 , w2483 );
and ( w2509 , w2507 , w2528 );
and ( w2510 , w2505 , w2509 );
not ( w2511 , w2499 );
and ( w2512 , w2511 , w2510 );
nor ( w2513 , w2506 , w1615 );
and ( w2514 , w2513 , w2528 );
and ( w2515 , w2512 , w2514 );
and ( w2516 , w2515 , w1624 );
and ( w2517 , w2516 , w1640 );
and ( w2518 , w2517 , w2514 );
not ( w2519 , w2492 );
and ( w2520 , w2519 , w2518 );
and ( w2521 , w1624 , w2520 );
not ( w2522 , w1821 );
and ( w2523 , w2522 , w2490 );
and ( w2524 , w1826 , w2540 );
and ( w2525 , w2521 , w2524 );
not ( w2526 , w2506 );
and ( w2527 , w2526 , w1623 );
not ( w2528 , w2508 );
and ( w2529 , w2527 , w2528 );
not ( w2530 , w2070 );
and ( w2531 , w2530 , w2489 );
not ( w2532 , w2531 );
and ( w2533 , w2529 , w2532 );
and ( w2534 , w2521 , w2533 );
and ( w2535 , w2534 , w2529 );
and ( w2536 , w2535 , w2521 );
and ( w2537 , w2540 , w2503 );
and ( w2538 , w2537 , w2509 );
and ( w2539 , w1869 , w2538 );
not ( w2540 , w2523 );
and ( w2541 , w2539 , w2540 );
and ( w2542 , w2536 , w2541 );
and ( w2543 , w2524 , w2529 );
and ( w2544 , w2542 , w2543 );
and ( w2545 , w2544 , w2529 );
and ( w2546 , w2541 , w2521 );
and ( w2547 , w2546 , w2533 );
and ( w2548 , w2545 , w2547 );
and ( w2549 , w2548 , w2521 );
and ( t_0 , w2525 , w2549 );
nor ( w2550 , w207 , g7 );
nor ( w2551 , g6 , g7 );
nor ( w2552 , w2551 , w52 );
and ( w2553 , w2552 , w11092 );
nor ( w2554 , w2553 , g5 );
and ( w2555 , w2554 , w12934 );
nor ( w2556 , w2555 , g5 );
and ( w2557 , w2556 , w12934 );
not ( w2558 , w2557 );
and ( w2559 , w2550 , w2558 );
nor ( w2560 , w2559 , g5 );
and ( w2561 , w2560 , w12934 );
not ( w2562 , w66 );
and ( w2563 , w1 , w2562 );
nor ( w2564 , w2563 , g3 );
and ( w2565 , w2564 , w6138 );
and ( w2566 , w2565 , w6144 );
nor ( w2567 , w2561 , w2566 );
not ( w2568 , w12 );
and ( w2569 , w2568 , g7 );
not ( w2570 , w2569 );
and ( w2571 , w2570 , w52 );
and ( w2572 , w2571 , w11092 );
nor ( w2573 , w2572 , w14 );
not ( w2574 , w2573 );
and ( w2575 , w2567 , w2574 );
nor ( w2576 , w8 , w14 );
nor ( w2577 , w212 , w2557 );
nor ( w2578 , w2577 , g5 );
and ( w2579 , w2578 , w12934 );
nor ( w2580 , w2576 , w2579 );
not ( w2581 , w2580 );
and ( w2582 , w2581 , w2573 );
nor ( w2583 , w8 , w1 );
and ( w2584 , w10 , w2583 );
nor ( w2585 , w212 , g5 );
and ( w2586 , w2585 , w12934 );
nor ( w2587 , w2584 , w2586 );
and ( w2588 , w5101 , w2587 );
nor ( w2589 , w2588 , w2575 );
and ( w2590 , w8 , w7419 );
and ( w2591 , w2554 , w2590 );
and ( w2592 , w2591 , w7419 );
and ( w2593 , w2589 , w6110 );
nor ( w2594 , w151 , g16 );
nor ( w2595 , w21 , g17 );
nor ( w2596 , w2594 , w2595 );
and ( w2597 , w2596 , w3811 );
and ( w2598 , g18 , w3811 );
and ( w2599 , w2598 , g19 );
nor ( w2600 , w2597 , w2599 );
and ( w2601 , w2600 , w8363 );
nor ( w2602 , w2601 , w31 );
nor ( w2603 , w2602 , w33 );
nor ( w2604 , w2603 , w37 );
nor ( w2605 , w2604 , w39 );
nor ( w2606 , w2605 , w31 );
nor ( w2607 , w2606 , w33 );
nor ( w2608 , w2607 , w37 );
nor ( w2609 , w2608 , w39 );
nor ( w2610 , w2609 , w41 );
nor ( w2611 , w2610 , w45 );
nor ( w2612 , w2611 , w48 );
and ( w2613 , w2612 , w12144 );
and ( w2614 , g10 , w13477 );
and ( w2615 , w11261 , g11 );
nor ( w2616 , w2614 , w2615 );
nor ( w2617 , w2613 , w2616 );
and ( w2618 , w2617 , w11166 );
nor ( w2619 , w485 , w2618 );
nor ( w2620 , w2619 , w19 );
and ( w2621 , w2727 , g5 );
not ( w2622 , w2621 );
and ( w2623 , w2622 , g5 );
nor ( w2624 , w2623 , w2553 );
and ( w2625 , w2620 , w2624 );
and ( w2626 , w2625 , w2587 );
nor ( w2627 , w2626 , w2575 );
and ( w2628 , w2627 , w6110 );
and ( w2629 , w4206 , g33 );
and ( w2630 , w2629 , g32 );
not ( w2631 , w2630 );
and ( w2632 , w2631 , g32 );
and ( w2633 , w2632 , g33 );
and ( w2634 , w8 , w11082 );
nor ( w2635 , w2634 , g2 );
not ( w2636 , g1 );
and ( w2637 , w2635 , w2636 );
and ( w2638 , w2641 , g5 );
nor ( w2639 , w2638 , w5 );
nor ( w2640 , w2639 , g7 );
not ( w2641 , w10 );
and ( w2642 , w2641 , g7 );
nor ( w2643 , w2640 , w2642 );
not ( w2644 , w2637 );
and ( w2645 , w2644 , w2643 );
not ( w2646 , w2645 );
and ( w2647 , w2646 , g32 );
not ( w2648 , w2647 );
and ( w2649 , w2648 , g32 );
and ( w2650 , w2633 , w5094 );
not ( w2651 , w2650 );
and ( w2652 , w2651 , w312 );
and ( w2653 , w2652 , w12717 );
and ( w2654 , w45 , w2587 );
nor ( w2655 , w8 , g3 );
and ( w2656 , w2655 , w6138 );
and ( w2657 , w2656 , w3175 );
nor ( w2658 , w8 , w2657 );
not ( w2659 , w2551 );
and ( w2660 , w8 , w2659 );
nor ( w2661 , w2660 , w14 );
not ( w2662 , w2661 );
and ( w2663 , w2658 , w2662 );
nor ( w2664 , w2663 , w2575 );
not ( w2665 , w2654 );
and ( w2666 , w2665 , w2664 );
nor ( w2667 , w274 , w2605 );
and ( w2668 , w2667 , w7485 );
and ( w2669 , w2668 , w12424 );
and ( w2670 , w2669 , w7803 );
nor ( w2671 , w2670 , w39 );
and ( w2672 , w11347 , w37 );
nor ( w2673 , w2672 , w41 );
and ( w2674 , w2673 , w3803 );
and ( w2675 , w2671 , w5422 );
and ( w2676 , w2675 , w12117 );
nor ( w2677 , w2676 , w43 );
not ( w2678 , w2677 );
and ( w2679 , w2678 , w2624 );
nor ( w2680 , w2679 , w2592 );
nor ( w2681 , w2666 , w2680 );
nor ( w2682 , w2681 , w2592 );
nor ( w2683 , w43 , w2682 );
nor ( w2684 , w2666 , w45 );
nor ( w2685 , w2684 , w2592 );
and ( w2686 , w2685 , w2582 );
and ( w2687 , w2686 , w2573 );
and ( w2688 , w2687 , w6110 );
not ( w2689 , w2683 );
and ( w2690 , w2689 , w2688 );
and ( w2691 , w2690 , w2582 );
not ( w2692 , w2691 );
and ( w2693 , w2692 , w2587 );
nor ( w2694 , w2693 , w2575 );
and ( w2695 , w2694 , w6110 );
nor ( w2696 , w2575 , w2592 );
and ( w2697 , w2695 , w2696 );
and ( w2698 , w2697 , w2666 );
and ( w2699 , w2698 , w12144 );
nor ( w2700 , w2699 , w2680 );
and ( w2701 , w2700 , w12144 );
nor ( w2702 , w2701 , w2592 );
and ( w2703 , w2702 , w2688 );
nor ( w2704 , w105 , w2703 );
and ( w2705 , w12921 , w2704 );
and ( w2706 , w8363 , w2705 );
not ( w2707 , w2706 );
and ( w2708 , w2707 , w2582 );
not ( w2709 , w2708 );
and ( w2710 , w2709 , w2624 );
and ( w2711 , w2710 , w2587 );
nor ( w2712 , w2711 , w2575 );
and ( w2713 , w2712 , w6110 );
and ( w2714 , w2713 , w19 );
not ( w2715 , w2714 );
and ( w2716 , w2715 , w310 );
and ( w2717 , w2716 , w312 );
and ( w2718 , w340 , w2741 );
and ( w2719 , w5101 , w2587 );
nor ( w2720 , w2719 , w2575 );
and ( w2721 , w2720 , w6110 );
not ( w2722 , w2718 );
and ( w2723 , w2722 , w2721 );
and ( w2724 , g34 , g35 );
nor ( w2725 , w69 , w2566 );
and ( w2726 , w2725 , g5 );
not ( w2727 , w69 );
and ( w2728 , w2727 , g7 );
nor ( w2729 , w2728 , w8 );
nor ( w2730 , w2729 , w2586 );
nor ( w2731 , w2551 , w2730 );
nor ( w2732 , w2731 , g5 );
and ( w2733 , w2732 , w2587 );
nor ( w2734 , w2726 , w2733 );
and ( w2735 , w2734 , w6003 );
nor ( w2736 , w2724 , w2735 );
and ( w2737 , w2736 , w2587 );
nor ( w2738 , w2737 , w2575 );
and ( w2739 , w2738 , w6110 );
nor ( w2740 , w2723 , w2739 );
not ( w2741 , w624 );
and ( w2742 , w340 , w2741 );
not ( w2743 , w2742 );
and ( w2744 , w2743 , w2721 );
nor ( w2745 , w2744 , w2739 );
and ( w2746 , w2745 , w5968 );
not ( w2747 , w2746 );
and ( w2748 , w2747 , w2582 );
not ( w2749 , w2748 );
and ( w2750 , w2749 , w2587 );
nor ( w2751 , w2750 , w2575 );
and ( w2752 , w2751 , w6110 );
not ( w2753 , w2740 );
and ( w2754 , w2753 , w2752 );
nor ( w2755 , w377 , w2573 );
and ( w2756 , w12921 , w2755 );
not ( w2757 , w2756 );
and ( w2758 , w2757 , w2573 );
and ( w2759 , w2754 , w2758 );
and ( w2760 , w2759 , w18 );
nor ( w2761 , w20 , w2760 );
and ( w2762 , w2761 , w5968 );
not ( w2763 , w2762 );
and ( w2764 , w2763 , w2582 );
not ( w2765 , w2764 );
and ( w2766 , w2765 , w2624 );
and ( w2767 , w2766 , w2587 );
nor ( w2768 , w2767 , w2575 );
and ( w2769 , w2768 , w6110 );
and ( w2770 , w2758 , w2664 );
and ( w2771 , w2770 , w2582 );
not ( w2772 , w2771 );
and ( w2773 , w2772 , w2587 );
nor ( w2774 , w2773 , w2575 );
and ( w2775 , w2774 , w6110 );
and ( w2776 , w2769 , w2775 );
and ( w2777 , w2776 , w18 );
and ( w2778 , w3811 , w272 );
and ( w2779 , g14 , g15 );
nor ( w2780 , w2779 , g17 );
nor ( w2781 , w2780 , w274 );
and ( w2782 , w2781 , g19 );
and ( w2783 , w2781 , w9197 );
nor ( w2784 , w2782 , w2783 );
nor ( w2785 , w2784 , w428 );
not ( w2786 , g16 );
and ( w2787 , w2786 , g17 );
nor ( w2788 , w2787 , w2780 );
and ( w2789 , w2788 , w11132 );
nor ( w2790 , w2789 , g19 );
and ( w2791 , w2790 , g18 );
not ( w2792 , w2791 );
and ( w2793 , w2792 , g18 );
not ( w2794 , w2789 );
and ( w2795 , w2794 , g19 );
not ( w2796 , w2795 );
and ( w2797 , w2796 , g19 );
nor ( w2798 , w2793 , w2797 );
and ( w2799 , w2798 , g20 );
nor ( w2800 , w2798 , w274 );
not ( w2801 , w2800 );
and ( w2802 , w2801 , g18 );
not ( w2803 , w2802 );
and ( w2804 , w2803 , g18 );
and ( w2805 , w2797 , w3811 );
not ( w2806 , w2805 );
and ( w2807 , w2806 , g19 );
not ( w2808 , w2807 );
and ( w2809 , w2808 , g19 );
nor ( w2810 , w2804 , w2809 );
nor ( w2811 , w2810 , w272 );
and ( w2812 , w3624 , g21 );
not ( w2813 , w2812 );
and ( w2814 , w2813 , g21 );
nor ( w2815 , w2814 , g20 );
nor ( w2816 , w2815 , w31 );
not ( w2817 , w2816 );
and ( w2818 , w2817 , w2587 );
nor ( w2819 , w2799 , w2818 );
and ( w2820 , w2819 , w3811 );
not ( w2821 , w2820 );
and ( w2822 , w2821 , g18 );
not ( w2823 , w2822 );
and ( w2824 , w2823 , g18 );
and ( w2825 , w2824 , w9197 );
nor ( w2826 , w2596 , g18 );
and ( w2827 , w2826 , w11347 );
and ( w2828 , w2827 , w8363 );
not ( w2829 , w2809 );
and ( w2830 , w2829 , w2828 );
nor ( w2831 , w2830 , w274 );
nor ( w2832 , w2831 , g18 );
and ( w2833 , w2832 , g19 );
nor ( w2834 , w2833 , g18 );
and ( w2835 , w2834 , g19 );
nor ( w2836 , w2835 , w2735 );
not ( w2837 , w2836 );
and ( w2838 , w2837 , w2582 );
not ( w2839 , w2838 );
and ( w2840 , w2839 , w2624 );
and ( w2841 , w2840 , w2587 );
nor ( w2842 , w2841 , w2575 );
and ( w2843 , w2842 , w6110 );
nor ( w2844 , w2825 , w2843 );
nor ( w2845 , w2844 , w272 );
and ( w2846 , w2845 , w7485 );
and ( w2847 , w2846 , w12424 );
nor ( w2848 , w2847 , w2735 );
not ( w2849 , w2848 );
and ( w2850 , w2849 , w2582 );
not ( w2851 , w2850 );
and ( w2852 , w2851 , w2624 );
and ( w2853 , w2852 , w2587 );
nor ( w2854 , w2853 , w2575 );
and ( w2855 , w2854 , w6110 );
and ( w2856 , w2785 , w2855 );
and ( w2857 , w2856 , w12085 );
and ( w2858 , w2857 , w7485 );
nor ( w2859 , w2858 , w2735 );
not ( w2860 , w2859 );
and ( w2861 , w2860 , w2582 );
not ( w2862 , w2861 );
and ( w2863 , w2862 , w2624 );
and ( w2864 , w2863 , w2587 );
nor ( w2865 , w2864 , w2575 );
and ( w2866 , w2865 , w6110 );
nor ( w2867 , w2778 , w2866 );
nor ( w2868 , w2867 , w35 );
and ( w2869 , w2868 , w7485 );
and ( w2870 , w2869 , w12424 );
and ( w2871 , w2870 , w7803 );
nor ( w2872 , w2871 , w39 );
and ( w2873 , w2872 , w5422 );
and ( w2874 , w2873 , w5370 );
nor ( w2875 , w2874 , w43 );
nor ( w2876 , w2875 , w2735 );
not ( w2877 , w2876 );
and ( w2878 , w2877 , w2582 );
not ( w2879 , w2878 );
and ( w2880 , w2879 , w2624 );
and ( w2881 , w2880 , w2587 );
nor ( w2882 , w2881 , w2575 );
and ( w2883 , w2882 , w6110 );
and ( w2884 , w2883 , w12142 );
nor ( w2885 , w2884 , w2735 );
and ( w2886 , w2885 , w2624 );
and ( w2887 , w2886 , w2587 );
nor ( w2888 , w2887 , w2575 );
nor ( w2889 , w105 , w2888 );
and ( w2890 , w2752 , w2664 );
and ( w2891 , w2890 , w2582 );
not ( w2892 , w2891 );
and ( w2893 , w2892 , w2587 );
nor ( w2894 , w2893 , w2575 );
and ( w2895 , w2894 , w6110 );
not ( w2896 , w2889 );
and ( w2897 , w2896 , w2895 );
nor ( w2898 , w2897 , w19 );
and ( w2899 , w2898 , w485 );
not ( w2900 , w2899 );
and ( w2901 , w2900 , w2713 );
and ( w2902 , w2901 , w6110 );
not ( w2903 , w2902 );
and ( w2904 , w310 , w2903 );
and ( w2905 , w2904 , w12532 );
and ( w2906 , g28 , w13333 );
nor ( w2907 , w2905 , w2906 );
nor ( w2908 , w134 , w2906 );
and ( w2909 , w2907 , w2908 );
not ( w2910 , w2909 );
and ( w2911 , w2910 , w377 );
and ( w2912 , w35 , w12424 );
and ( w2913 , w2912 , w7803 );
and ( w2914 , w11140 , w2913 );
not ( w2915 , w2914 );
and ( w2916 , w2915 , w2666 );
nor ( w2917 , w2916 , w2674 );
and ( w2918 , w2917 , w12117 );
and ( w2919 , w2918 , w12144 );
nor ( w2920 , w2919 , w2592 );
and ( w2921 , w2920 , w2573 );
and ( w2922 , w2921 , w6110 );
and ( w2923 , w2695 , w2922 );
and ( w2924 , w2923 , w2582 );
not ( w2925 , w2924 );
and ( w2926 , w2925 , w2587 );
nor ( w2927 , w2926 , w2575 );
and ( w2928 , w2927 , w6110 );
and ( w2929 , w2928 , w2922 );
and ( w2930 , w2929 , w2688 );
and ( w2931 , w2930 , w6110 );
nor ( w2932 , w20 , w2931 );
not ( w2933 , w2932 );
and ( w2934 , w2933 , w2582 );
not ( w2935 , w2934 );
and ( w2936 , w2935 , w2624 );
and ( w2937 , w2936 , w2587 );
nor ( w2938 , w2937 , w2575 );
and ( w2939 , w2938 , w6110 );
and ( w2940 , w2695 , w2939 );
and ( w2941 , w2940 , w2666 );
nor ( w2942 , w2941 , w2680 );
not ( w2943 , w2942 );
and ( w2944 , w2943 , w2688 );
and ( w2945 , w2944 , w2775 );
nor ( w2946 , w43 , w2945 );
nor ( w2947 , w2946 , w2592 );
and ( w2948 , w2947 , w11166 );
and ( w2949 , w2948 , w12498 );
and ( w2950 , w2758 , w12921 );
and ( w2951 , w2950 , w105 );
not ( w2952 , w2951 );
and ( w2953 , w2952 , g13 );
not ( w2954 , w2953 );
and ( w2955 , w2954 , w105 );
and ( w2956 , w2955 , g13 );
not ( w2957 , w2956 );
and ( w2958 , w2957 , w2624 );
not ( w2959 , w2958 );
and ( w2960 , w2959 , w2573 );
and ( w2961 , w2960 , w6110 );
nor ( w2962 , w2949 , w2961 );
and ( w2963 , w2962 , w12498 );
and ( w2964 , w12921 , w2963 );
not ( w2965 , w2964 );
and ( w2966 , w2965 , w2582 );
not ( w2967 , w2966 );
and ( w2968 , w2967 , w2624 );
and ( w2969 , w2968 , w2587 );
nor ( w2970 , w2969 , w2575 );
and ( w2971 , w2970 , w6110 );
not ( w2972 , w2911 );
and ( w2973 , w2972 , w2971 );
and ( w2974 , w18 , w2587 );
not ( w2975 , w2974 );
and ( w2976 , w2975 , w2664 );
and ( w2977 , w2973 , w2976 );
nor ( w2978 , w20 , w2977 );
and ( w2979 , w8363 , w2978 );
and ( w2980 , w2979 , w239 );
and ( w2981 , w2950 , w18 );
nor ( w2982 , w2981 , w20 );
not ( w2983 , w2982 );
and ( w2984 , w2983 , w18 );
and ( w2985 , w2984 , w12921 );
and ( w2986 , w18 , w12921 );
nor ( w2987 , w2986 , w2735 );
not ( w2988 , w2987 );
and ( w2989 , w2988 , w2582 );
not ( w2990 , w2989 );
and ( w2991 , w2990 , w2624 );
and ( w2992 , w2991 , w2587 );
nor ( w2993 , w2992 , w2575 );
and ( w2994 , w2993 , w6110 );
and ( w2995 , w2985 , w2994 );
and ( w2996 , w12144 , w2681 );
not ( w2997 , w2996 );
and ( w2998 , w2997 , w2688 );
nor ( w2999 , w20 , w2998 );
not ( w3000 , w2999 );
and ( w3001 , w3000 , w2582 );
not ( w3002 , w3001 );
and ( w3003 , w3002 , w2624 );
and ( w3004 , w3003 , w2587 );
nor ( w3005 , w3004 , w2575 );
and ( w3006 , w2770 , w3005 );
and ( w3007 , w3006 , w2976 );
nor ( w3008 , w3007 , w20 );
nor ( w3009 , w3008 , w105 );
nor ( w3010 , w3009 , w2961 );
and ( w3011 , w3010 , w5968 );
not ( w3012 , w3011 );
and ( w3013 , w3012 , w2582 );
not ( w3014 , w3013 );
and ( w3015 , w3014 , w2587 );
nor ( w3016 , w3015 , w2575 );
and ( w3017 , w3016 , w6110 );
and ( w3018 , w3017 , w11166 );
nor ( w3019 , w3018 , w2961 );
not ( w3020 , w3019 );
and ( w3021 , w3020 , w2582 );
not ( w3022 , w3021 );
and ( w3023 , w3022 , w2624 );
and ( w3024 , w3023 , w2587 );
nor ( w3025 , w3024 , w2575 );
and ( w3026 , w3025 , w6110 );
nor ( w3027 , w2995 , w3026 );
and ( w3028 , w20 , w11166 );
and ( w3029 , w2890 , w3005 );
and ( w3030 , w2752 , w2664 );
and ( w3031 , w3030 , w3005 );
and ( w3032 , w3031 , w2976 );
nor ( w3033 , w3032 , w20 );
not ( w3034 , w3033 );
and ( w3035 , w3034 , w3026 );
nor ( w3036 , w3035 , w2735 );
not ( w3037 , w3036 );
and ( w3038 , w3037 , w2582 );
not ( w3039 , w3038 );
and ( w3040 , w3039 , w2587 );
nor ( w3041 , w3040 , w2575 );
and ( w3042 , w3041 , w6110 );
and ( w3043 , w3029 , w3042 );
not ( w3044 , w2754 );
and ( w3045 , w105 , w3044 );
not ( w3046 , w3045 );
and ( w3047 , w3046 , w2976 );
and ( w3048 , w3047 , w3026 );
nor ( w3049 , w3048 , w20 );
and ( w3050 , w3049 , w5968 );
not ( w3051 , w3050 );
and ( w3052 , w3051 , w2582 );
not ( w3053 , w3052 );
and ( w3054 , w3053 , w2624 );
and ( w3055 , w3054 , w2587 );
nor ( w3056 , w3055 , w2575 );
and ( w3057 , w3056 , w6110 );
and ( w3058 , w3043 , w3057 );
and ( w3059 , w3058 , w3026 );
nor ( w3060 , w3059 , w2769 );
and ( w3061 , w3060 , w5968 );
not ( w3062 , w3061 );
and ( w3063 , w3062 , w2582 );
not ( w3064 , w3063 );
and ( w3065 , w3064 , w2587 );
nor ( w3066 , w3065 , w2575 );
and ( w3067 , w3066 , w6110 );
not ( w3068 , w3028 );
and ( w3069 , w3068 , w3067 );
and ( w3070 , w3042 , w11166 );
and ( w3071 , w3070 , w8640 );
not ( w3072 , w3071 );
and ( w3073 , w3072 , w377 );
not ( w3074 , w3073 );
and ( w3075 , w3074 , w3026 );
nor ( w3076 , w3075 , w2735 );
not ( w3077 , w3076 );
and ( w3078 , w3077 , w2582 );
not ( w3079 , w3078 );
and ( w3080 , w3079 , w2624 );
and ( w3081 , w3080 , w2587 );
nor ( w3082 , w3081 , w2575 );
and ( w3083 , w3082 , w6110 );
nor ( w3084 , w3069 , w3083 );
nor ( w3085 , w3084 , w2592 );
not ( w3086 , w3085 );
and ( w3087 , w3086 , g31 );
and ( w3088 , w310 , w3087 );
and ( w3089 , w3005 , w2976 );
nor ( w3090 , w20 , w2573 );
not ( w3091 , w3090 );
and ( w3092 , w3091 , w2582 );
not ( w3093 , w3092 );
and ( w3094 , w3093 , w2624 );
not ( w3095 , w3094 );
and ( w3096 , w3095 , w2573 );
and ( w3097 , w3096 , w6110 );
and ( w3098 , w3097 , w2664 );
nor ( w3099 , w20 , w3098 );
not ( w3100 , w3099 );
and ( w3101 , w3100 , w2582 );
not ( w3102 , w3101 );
and ( w3103 , w3102 , w2624 );
and ( w3104 , w3103 , w2587 );
nor ( w3105 , w3104 , w2575 );
and ( w3106 , w3105 , w6110 );
and ( w3107 , w3089 , w3106 );
and ( w3108 , w2573 , w18 );
nor ( w3109 , w20 , w3108 );
and ( w3110 , w3109 , w2624 );
not ( w3111 , w3110 );
and ( w3112 , w3111 , w2573 );
and ( w3113 , w3112 , w6110 );
and ( w3114 , w3113 , w18 );
and ( w3115 , w3114 , w2573 );
and ( w3116 , w3115 , w6110 );
nor ( w3117 , w3107 , w3116 );
nor ( w3118 , w3117 , w105 );
nor ( w3119 , w3118 , w2961 );
not ( w3120 , w3119 );
and ( w3121 , w3120 , w2582 );
not ( w3122 , w3121 );
and ( w3123 , w3122 , w2587 );
nor ( w3124 , w3123 , w2575 );
and ( w3125 , w3124 , w11166 );
nor ( w3126 , w3125 , w2961 );
not ( w3127 , w3126 );
and ( w3128 , w3127 , w2582 );
not ( w3129 , w3128 );
and ( w3130 , w3129 , w2587 );
nor ( w3131 , w3130 , w2575 );
not ( w3132 , w3088 );
and ( w3133 , w3132 , w3131 );
nor ( w3134 , w3133 , w308 );
and ( w3135 , w3134 , w11852 );
and ( w3136 , w3135 , w12037 );
and ( w3137 , w3136 , w5968 );
not ( w3138 , w3137 );
and ( w3139 , w3138 , w2582 );
not ( w3140 , w3139 );
and ( w3141 , w3140 , w2624 );
and ( w3142 , w3141 , w2587 );
nor ( w3143 , w3142 , w2575 );
and ( w3144 , w3143 , w6110 );
not ( w3145 , w3027 );
and ( w3146 , w3145 , w3144 );
and ( w3147 , w310 , w8848 );
and ( w3148 , w3147 , g32 );
and ( w3149 , w3148 , g33 );
nor ( w3150 , w19 , w312 );
and ( w3151 , w3150 , w2587 );
nor ( w3152 , w3149 , w3151 );
nor ( w3153 , w3152 , w105 );
and ( w3154 , w3153 , w2587 );
and ( w3155 , w3154 , w377 );
and ( w3156 , w3155 , w12080 );
and ( w3157 , w377 , w3156 );
nor ( w3158 , w384 , w19 );
and ( w3159 , w789 , w13333 );
not ( w3160 , w3159 );
and ( w3161 , g28 , w3160 );
nor ( w3162 , w3161 , w377 );
and ( w3163 , w3162 , w12080 );
and ( w3164 , w3163 , w20 );
and ( w3165 , w3162 , g10 );
and ( w3166 , w67 , w3175 );
nor ( w3167 , w3166 , w8 );
nor ( w3168 , w208 , g7 );
nor ( w3169 , w3168 , g7 );
nor ( w3170 , w3167 , w3169 );
and ( w3171 , w3170 , w7419 );
nor ( w3172 , w3171 , w2592 );
nor ( w3173 , w66 , w3169 );
and ( w3174 , w3173 , w2643 );
not ( w3175 , w1 );
and ( w3176 , w3174 , w3175 );
and ( w3177 , w3176 , w10 );
nor ( w3178 , w2609 , w48 );
nor ( w3179 , w20 , w3178 );
and ( w3180 , w3179 , w2624 );
nor ( w3181 , w3180 , w41 );
nor ( w3182 , w3181 , w45 );
nor ( w3183 , w3182 , w43 );
not ( w3184 , w3177 );
and ( w3185 , w3184 , w3183 );
and ( w3186 , w3185 , w11166 );
and ( w3187 , w3172 , w3186 );
and ( w3188 , w3187 , w12142 );
not ( w3189 , w3188 );
and ( w3190 , w3189 , w3162 );
and ( w3191 , w3190 , w12717 );
and ( w3192 , w3191 , w12919 );
and ( w3193 , w3192 , w13477 );
and ( w3194 , w3193 , g33 );
and ( w3195 , w3194 , w11166 );
and ( w3196 , w3195 , w789 );
and ( w3197 , w3196 , w11261 );
and ( w3198 , w3197 , w13477 );
and ( w3199 , w3198 , w12080 );
and ( w3200 , w3199 , w13477 );
and ( w3201 , w3200 , g33 );
and ( w3202 , w3201 , w11166 );
and ( w3203 , w3202 , w12717 );
and ( w3204 , w3203 , w11261 );
and ( w3205 , w3204 , w2587 );
and ( w3206 , w3205 , w13477 );
nor ( w3207 , w3165 , w3206 );
nor ( w3208 , w3207 , g11 );
and ( w3209 , w3208 , w12717 );
and ( w3210 , w3209 , w12080 );
and ( w3211 , w3210 , g33 );
and ( w3212 , w3211 , w12498 );
and ( w3213 , w3212 , w2587 );
not ( w3214 , w3213 );
and ( w3215 , w3214 , w2664 );
and ( w3216 , w3215 , w13477 );
not ( w3217 , w3216 );
and ( w3218 , w3163 , w3217 );
and ( w3219 , w12498 , w3218 );
and ( w3220 , w3219 , g33 );
and ( w3221 , w3220 , w12717 );
and ( w3222 , w3221 , w12080 );
nor ( w3223 , w2673 , w39 );
nor ( w3224 , w43 , w3223 );
not ( w3225 , w3224 );
and ( w3226 , w3222 , w3225 );
and ( w3227 , w3226 , w12117 );
and ( w3228 , w3227 , w43 );
and ( w3229 , w12142 , w2587 );
not ( w3230 , w3229 );
and ( w3231 , w3230 , w2664 );
nor ( w3232 , w39 , w3231 );
nor ( w3233 , w3232 , w2592 );
and ( w3234 , w3163 , w5366 );
and ( w3235 , w3234 , w3833 );
and ( w3236 , w3235 , w12498 );
not ( w3237 , w3236 );
and ( w3238 , w3237 , w2573 );
not ( w3239 , w3238 );
and ( w3240 , w3162 , w3239 );
and ( w3241 , w3215 , w12921 );
and ( w3242 , w3241 , w11261 );
and ( w3243 , w3242 , w13477 );
nor ( w3244 , w3206 , w20 );
not ( w3245 , w3206 );
and ( w3246 , w2950 , w3245 );
and ( w3247 , w3246 , w12921 );
and ( w3248 , w3247 , w105 );
not ( w3249 , w3248 );
and ( w3250 , w3249 , g13 );
not ( w3251 , w3250 );
and ( w3252 , w3251 , w105 );
and ( w3253 , w3252 , g13 );
nor ( w3254 , w377 , w3253 );
and ( w3255 , w3254 , w2624 );
not ( w3256 , w3255 );
and ( w3257 , w3256 , w2573 );
and ( w3258 , w3257 , w6110 );
nor ( w3259 , w3244 , w3258 );
nor ( w3260 , w3259 , g10 );
and ( w3261 , w3260 , w13477 );
nor ( w3262 , w377 , w3261 );
not ( w3263 , w3262 );
and ( w3264 , w3263 , w2573 );
and ( w3265 , w3264 , w6110 );
nor ( w3266 , w3243 , w3265 );
and ( w3267 , w12498 , w3266 );
not ( w3268 , w3267 );
and ( w3269 , w3268 , w2573 );
and ( w3270 , w3269 , w6110 );
nor ( w3271 , w3270 , w3231 );
nor ( w3272 , w3271 , w48 );
not ( w3273 , w3272 );
and ( w3274 , w3273 , g33 );
and ( w3275 , w3274 , w12717 );
and ( w3276 , w3275 , w12080 );
and ( w3277 , w3240 , w3276 );
and ( w3278 , w3277 , w5366 );
and ( w3279 , w3278 , w5422 );
and ( w3280 , w3279 , w11140 );
and ( w3281 , w3280 , w12117 );
and ( w3282 , w3162 , w11261 );
and ( w3283 , w3282 , g11 );
not ( w3284 , w3283 );
and ( w3285 , w3284 , w3215 );
nor ( w3286 , w3285 , g9 );
not ( w3287 , g8 );
and ( w3288 , w3286 , w3287 );
and ( w3289 , w3288 , w48 );
and ( w3290 , w3289 , w12717 );
and ( w3291 , w3290 , w12080 );
and ( w3292 , w3291 , w12919 );
and ( w3293 , w3292 , g33 );
and ( w3294 , w3293 , w12498 );
and ( w3295 , w3294 , w2587 );
not ( w3296 , w3295 );
and ( w3297 , w3296 , w2664 );
not ( w3298 , w3281 );
and ( w3299 , w3298 , w3297 );
and ( w3300 , w3299 , w8848 );
and ( w3301 , w3300 , w11166 );
and ( w3302 , w3301 , w12921 );
nor ( w3303 , w377 , w3302 );
and ( w3304 , w3303 , g33 );
and ( w3305 , w3304 , w12717 );
and ( w3306 , w3305 , w12080 );
not ( w3307 , w3306 );
and ( w3308 , w3307 , w2573 );
and ( w3309 , w3308 , w6110 );
nor ( w3310 , w2605 , w37 );
nor ( w3311 , w3310 , w3231 );
not ( w3312 , w3311 );
and ( w3313 , w3312 , w2573 );
and ( w3314 , w3313 , w12144 );
nor ( w3315 , w20 , w3314 );
and ( w3316 , w12498 , w3315 );
and ( w3317 , w3316 , w2624 );
not ( w3318 , w3317 );
and ( w3319 , w3318 , w2573 );
and ( w3320 , w3319 , w6110 );
and ( w3321 , w7803 , w3320 );
and ( w3322 , w3665 , w2587 );
nor ( w3323 , w48 , w3322 );
nor ( w3324 , w3323 , w20 );
and ( w3325 , w3321 , w3829 );
and ( w3326 , w3325 , w11166 );
nor ( w3327 , w20 , w3326 );
not ( w3328 , w3327 );
and ( w3329 , w3328 , w2573 );
and ( w3330 , w3329 , w6110 );
nor ( w3331 , w3309 , w3330 );
and ( w3332 , w3331 , w5366 );
and ( w3333 , w3332 , w5422 );
and ( w3334 , w3333 , w11140 );
and ( w3335 , w3334 , w12117 );
and ( w3336 , w3335 , w3833 );
not ( w3337 , w3336 );
and ( w3338 , w3337 , w3297 );
and ( w3339 , w3338 , w8848 );
and ( w3340 , w3339 , w11166 );
and ( w3341 , w3340 , w2976 );
nor ( w3342 , w20 , w3341 );
and ( w3343 , w12498 , w3342 );
and ( w3344 , w3343 , g33 );
and ( w3345 , w3344 , w12717 );
and ( w3346 , w3345 , w12080 );
and ( w3347 , w3346 , w2624 );
not ( w3348 , w3347 );
and ( w3349 , w3348 , w2573 );
and ( w3350 , w3349 , w6110 );
not ( w3351 , w3228 );
and ( w3352 , w3351 , w3350 );
and ( w3353 , w3350 , w2573 );
and ( w3354 , w3353 , w2976 );
nor ( w3355 , w20 , w3354 );
nor ( w3356 , w3355 , w105 );
nor ( w3357 , w377 , w3356 );
and ( w3358 , w3357 , w12080 );
and ( w3359 , w3358 , w2624 );
not ( w3360 , w3359 );
and ( w3361 , w3360 , w2573 );
and ( w3362 , w3361 , w6110 );
and ( w3363 , w3352 , w3362 );
not ( w3364 , w3363 );
and ( w3365 , w3364 , w3276 );
and ( w3366 , w3365 , w5597 );
and ( w3367 , w3366 , w12921 );
nor ( w3368 , w3367 , w105 );
nor ( w3369 , w377 , w3368 );
and ( w3370 , w12717 , w3369 );
and ( w3371 , w3370 , w12080 );
not ( w3372 , w3371 );
and ( w3373 , w3372 , w2573 );
and ( w3374 , w3373 , w6110 );
not ( w3375 , w3374 );
and ( w3376 , w3375 , w43 );
not ( w3377 , w3376 );
and ( w3378 , w3377 , w3350 );
not ( w3379 , w3378 );
and ( w3380 , w3379 , w3322 );
and ( w3381 , w3380 , w3833 );
and ( w3382 , w3381 , w5597 );
not ( w3383 , w3382 );
and ( w3384 , w3383 , w3297 );
nor ( w3385 , w20 , w3384 );
nor ( w3386 , w3362 , w3116 );
and ( w3387 , w12921 , w3386 );
and ( w3388 , w3387 , w3947 );
and ( w3389 , w12498 , w3388 );
and ( w3390 , w12717 , w3389 );
not ( w3391 , w3390 );
and ( w3392 , w3391 , w2573 );
and ( w3393 , w3392 , w11166 );
nor ( w3394 , w3393 , w2961 );
not ( w3395 , w3394 );
and ( w3396 , w3395 , w2573 );
not ( w3397 , w3385 );
and ( w3398 , w3397 , w3396 );
and ( w3399 , w3398 , w8848 );
and ( w3400 , w3399 , w11166 );
nor ( w3401 , w3400 , w2961 );
and ( w3402 , w12498 , w3401 );
and ( w3403 , w3402 , g33 );
and ( w3404 , w12717 , w3403 );
and ( w3405 , w3404 , w12080 );
not ( w3406 , w3405 );
and ( w3407 , w3406 , w2573 );
and ( w3408 , w3407 , w6110 );
not ( w3409 , w3164 );
and ( w3410 , w3409 , w3408 );
nor ( w3411 , w3410 , w2961 );
and ( w3412 , w3411 , w12498 );
and ( w3413 , w3412 , g33 );
and ( w3414 , w3413 , w12717 );
and ( w3415 , w3414 , w12080 );
not ( w3416 , w3415 );
and ( w3417 , w3416 , w2573 );
nor ( w3418 , w3417 , w19 );
nor ( w3419 , w20 , w2573 );
and ( w3420 , w19 , w3419 );
not ( w3421 , w3420 );
and ( w3422 , w3421 , w2582 );
not ( w3423 , w3422 );
and ( w3424 , w3423 , w2624 );
not ( w3425 , w3424 );
and ( w3426 , w3425 , w2573 );
and ( w3427 , w3426 , w6110 );
not ( w3428 , w3418 );
and ( w3429 , w3428 , w3427 );
and ( w3430 , w11852 , g29 );
and ( w3431 , w3430 , g28 );
and ( w3432 , w12717 , w3431 );
and ( w3433 , w3432 , w2587 );
and ( w3434 , w3429 , w3445 );
and ( w3435 , w3434 , w11852 );
nor ( w3436 , w3435 , w2735 );
not ( w3437 , w3436 );
and ( w3438 , w3437 , w2582 );
not ( w3439 , w3438 );
and ( w3440 , w3439 , w2587 );
nor ( w3441 , w3440 , w2575 );
and ( w3442 , w3441 , w12717 );
and ( w3443 , w3442 , w12498 );
and ( w3444 , w12717 , g31 );
not ( w3445 , w3433 );
and ( w3446 , w3444 , w3445 );
not ( w3447 , w3446 );
and ( w3448 , w3447 , w2587 );
and ( w3449 , w3448 , g30 );
and ( w3450 , w3449 , g31 );
and ( w3451 , w310 , w3450 );
and ( w3452 , g30 , w13206 );
not ( w3453 , w3452 );
and ( w3454 , w3453 , g30 );
and ( w3455 , w3454 , w13206 );
and ( w3456 , w12199 , g31 );
nor ( w3457 , w3456 , g30 );
and ( w3458 , w3457 , g31 );
nor ( w3459 , w3455 , w3458 );
and ( w3460 , w3459 , w13333 );
not ( w3461 , w3460 );
and ( w3462 , w3461 , w3417 );
nor ( w3463 , w3462 , w19 );
not ( w3464 , w3463 );
and ( w3465 , w3464 , w3427 );
nor ( w3466 , w3465 , w310 );
nor ( w3467 , w3466 , w3433 );
and ( w3468 , w3467 , w11852 );
nor ( w3469 , w3468 , w2735 );
not ( w3470 , w3469 );
and ( w3471 , w3470 , w2582 );
not ( w3472 , w3471 );
and ( w3473 , w3472 , w2587 );
nor ( w3474 , w3473 , w2575 );
not ( w3475 , w3451 );
and ( w3476 , w3475 , w3474 );
nor ( w3477 , w3476 , w2735 );
and ( w3478 , w3477 , w2587 );
nor ( w3479 , w3478 , w2575 );
nor ( w3480 , w3479 , w2735 );
and ( w3481 , w3480 , w2587 );
nor ( w3482 , w3481 , w2575 );
nor ( w3483 , w3443 , w3482 );
and ( w3484 , w3483 , w5968 );
and ( w3485 , w3484 , w2587 );
nor ( w3486 , w3485 , w2575 );
and ( w3487 , w3158 , w4464 );
and ( w3488 , w3417 , w12080 );
and ( w3489 , w3488 , w12498 );
nor ( w3490 , w3489 , w2735 );
and ( w3491 , w3490 , w2587 );
nor ( w3492 , w3491 , w2575 );
nor ( w3493 , w3482 , w3492 );
and ( w3494 , w12498 , w3097 );
and ( w3495 , w2908 , w377 );
and ( w3496 , w3495 , w13333 );
nor ( w3497 , w3496 , w2735 );
and ( w3498 , w3497 , w2587 );
nor ( w3499 , w3498 , w2575 );
and ( w3500 , w3499 , w6110 );
nor ( w3501 , w3494 , w3500 );
and ( w3502 , w384 , w3501 );
and ( w3503 , w3427 , w2582 );
not ( w3504 , w3503 );
and ( w3505 , w3504 , w2587 );
nor ( w3506 , w3505 , w2575 );
not ( w3507 , w3502 );
and ( w3508 , w3507 , w3506 );
nor ( w3509 , w3508 , w2735 );
not ( w3510 , w3509 );
and ( w3511 , w3510 , w2582 );
not ( w3512 , w3511 );
and ( w3513 , w3512 , w2587 );
nor ( w3514 , w3513 , w2575 );
and ( w3515 , w3514 , w6110 );
and ( w3516 , w3515 , w8640 );
and ( w3517 , w3516 , w19 );
and ( w3518 , w3517 , w2582 );
not ( w3519 , w3518 );
and ( w3520 , w3519 , w2624 );
and ( w3521 , w3520 , w2587 );
nor ( w3522 , w3521 , w2575 );
not ( w3523 , w3522 );
and ( w3524 , w3493 , w3523 );
not ( w3525 , w3517 );
and ( w3526 , w3525 , g11 );
not ( w3527 , w3526 );
and ( w3528 , w3527 , w19 );
and ( w3529 , w3528 , g11 );
nor ( w3530 , w3529 , w2735 );
not ( w3531 , w3530 );
and ( w3532 , w3531 , w2582 );
not ( w3533 , w3532 );
and ( w3534 , w3533 , w2624 );
and ( w3535 , w3534 , w2587 );
nor ( w3536 , w3535 , w2575 );
not ( w3537 , w3536 );
and ( w3538 , w3524 , w3537 );
and ( w3539 , w3538 , w12199 );
nor ( w3540 , w3539 , g30 );
nor ( w3541 , w3540 , g31 );
not ( w3542 , w3541 );
and ( w3543 , w3542 , w384 );
and ( w3544 , w3543 , w13206 );
not ( w3545 , w3474 );
and ( w3546 , w377 , w3545 );
not ( w3547 , w3546 );
and ( w3548 , w3547 , w3441 );
nor ( w3549 , w3548 , w19 );
not ( w3550 , w3549 );
and ( w3551 , w3550 , w3506 );
and ( w3552 , w3551 , w11852 );
nor ( w3553 , w3552 , w2735 );
not ( w3554 , w3553 );
and ( w3555 , w3554 , w2582 );
not ( w3556 , w3555 );
and ( w3557 , w3556 , w2587 );
nor ( w3558 , w3557 , w2575 );
nor ( w3559 , w3558 , w19 );
not ( w3560 , w3559 );
and ( w3561 , w3560 , w3506 );
and ( w3562 , w3561 , w11852 );
and ( w3563 , w3562 , w2647 );
not ( w3564 , w3563 );
and ( w3565 , w3564 , g32 );
not ( w3566 , w3565 );
and ( w3567 , w3566 , g32 );
and ( w3568 , w3567 , g33 );
nor ( w3569 , w3568 , w2735 );
not ( w3570 , w3569 );
and ( w3571 , w3570 , w2582 );
not ( w3572 , w3571 );
and ( w3573 , w3572 , w2624 );
and ( w3574 , w3573 , w2587 );
nor ( w3575 , w3574 , w2575 );
nor ( w3576 , w3544 , w3575 );
nor ( w3577 , w308 , w312 );
nor ( w3578 , g33 , w3577 );
not ( w3579 , w3578 );
and ( w3580 , w3579 , w2647 );
not ( w3581 , w2590 );
and ( w3582 , w3580 , w3581 );
not ( w3583 , w3576 );
and ( w3584 , w3583 , w3582 );
and ( w3585 , w3584 , w2647 );
not ( w3586 , w3585 );
and ( w3587 , w3586 , g32 );
not ( w3588 , w3587 );
and ( w3589 , w3588 , g32 );
and ( w3590 , w3589 , g33 );
nor ( w3591 , w3590 , w2735 );
not ( w3592 , w3591 );
and ( w3593 , w3592 , w2582 );
not ( w3594 , w3593 );
and ( w3595 , w3594 , w2624 );
and ( w3596 , w3595 , w2587 );
nor ( w3597 , w3596 , w2575 );
and ( w3598 , w384 , w3597 );
nor ( w3599 , w3598 , w3575 );
not ( w3600 , w3599 );
and ( w3601 , w3600 , w2582 );
not ( w3602 , w3601 );
and ( w3603 , w3602 , w2587 );
nor ( w3604 , w3603 , w2575 );
and ( w3605 , w3604 , w6110 );
not ( w3606 , w3487 );
and ( w3607 , w3606 , w3605 );
not ( w3608 , w3607 );
and ( w3609 , w3608 , g32 );
and ( w3610 , w3609 , g33 );
nor ( w3611 , w3610 , w2649 );
and ( w3612 , w2589 , w2582 );
not ( w3613 , w3612 );
and ( w3614 , w3613 , w2587 );
nor ( w3615 , w3614 , w2575 );
and ( w3616 , w19 , w3615 );
not ( w3617 , w3616 );
and ( w3618 , w3617 , g31 );
and ( w3619 , w3618 , w11852 );
and ( w3620 , w3619 , w310 );
nor ( w3621 , w255 , w19 );
not ( w3622 , w3621 );
and ( w3623 , w3622 , w2587 );
not ( w3624 , w2811 );
and ( w3625 , w3624 , g20 );
nor ( w3626 , w3625 , w2818 );
and ( w3627 , w3626 , w2922 );
and ( w3628 , w3627 , w7485 );
and ( w3629 , w3628 , w12424 );
nor ( w3630 , w3629 , w2735 );
not ( w3631 , w3630 );
and ( w3632 , w3631 , w2582 );
not ( w3633 , w3632 );
and ( w3634 , w3633 , w2624 );
and ( w3635 , w3634 , w2587 );
nor ( w3636 , w3635 , w2575 );
and ( w3637 , w3636 , w6110 );
and ( w3638 , w3637 , w7485 );
and ( w3639 , w3638 , w12424 );
nor ( w3640 , w3639 , w2735 );
and ( w3641 , w3640 , w2587 );
nor ( w3642 , w3641 , w2575 );
and ( w3643 , w3642 , w6110 );
and ( w3644 , w3637 , w3643 );
and ( w3645 , w3644 , w7485 );
and ( w3646 , w3645 , w12424 );
and ( w3647 , w3646 , w7803 );
nor ( w3648 , w3647 , w39 );
and ( w3649 , w3648 , w5370 );
not ( w3650 , w3649 );
and ( w3651 , w3650 , w2976 );
nor ( w3652 , w3651 , w3113 );
nor ( w3653 , w3652 , w2592 );
and ( w3654 , w3653 , w12921 );
and ( w3655 , w3654 , w8640 );
and ( w3656 , w3655 , w12144 );
and ( w3657 , w3656 , w12142 );
and ( w3658 , w3657 , w3106 );
and ( w3659 , w12921 , w3658 );
and ( w3660 , w3626 , w7485 );
and ( w3661 , w3660 , w12424 );
nor ( w3662 , w3661 , w39 );
nor ( w3663 , w3662 , w41 );
nor ( w3664 , w3663 , w2674 );
not ( w3665 , w3186 );
and ( w3666 , w3664 , w3665 );
not ( w3667 , w3666 );
and ( w3668 , w3667 , w2664 );
and ( w3669 , w3668 , w11261 );
and ( w3670 , w3669 , w13477 );
nor ( w3671 , w3670 , w48 );
nor ( w3672 , w3671 , w2592 );
and ( w3673 , w3672 , w12144 );
and ( w3674 , w3673 , w12142 );
nor ( w3675 , w3674 , w2961 );
and ( w3676 , w3675 , w5968 );
not ( w3677 , w3676 );
and ( w3678 , w3677 , w2582 );
not ( w3679 , w3678 );
and ( w3680 , w3679 , w2624 );
and ( w3681 , w3680 , w2587 );
nor ( w3682 , w3681 , w2575 );
and ( w3683 , w3682 , w6110 );
nor ( w3684 , w3683 , w3116 );
and ( w3685 , w12921 , w3684 );
and ( w3686 , w3685 , w5968 );
and ( w3687 , w3686 , w2624 );
and ( w3688 , w3687 , w2587 );
nor ( w3689 , w3688 , w2575 );
and ( w3690 , w12921 , w3689 );
and ( w3691 , w3690 , w12498 );
nor ( w3692 , w3691 , w2961 );
and ( w3693 , w3692 , w12498 );
and ( w3694 , w3693 , w5968 );
and ( w3695 , w3694 , w2587 );
nor ( w3696 , w3695 , w2575 );
nor ( w3697 , w3659 , w3696 );
nor ( w3698 , w3697 , w105 );
nor ( w3699 , w3698 , w2961 );
and ( w3700 , w3699 , w5968 );
and ( w3701 , w3700 , w2624 );
and ( w3702 , w3701 , w2587 );
nor ( w3703 , w3702 , w2575 );
and ( w3704 , w3703 , w6110 );
not ( w3705 , w3704 );
and ( w3706 , w3623 , w3705 );
and ( w3707 , w3706 , w255 );
and ( w3708 , w8848 , w3707 );
not ( w3709 , w3708 );
and ( w3710 , w3709 , w3615 );
nor ( w3711 , w3710 , w377 );
and ( w3712 , w3711 , w12717 );
and ( w3713 , w3712 , w11852 );
and ( w3714 , w3713 , w12037 );
and ( w3715 , w3714 , w5898 );
and ( w3716 , w3715 , w11166 );
and ( w3717 , w3716 , w5968 );
not ( w3718 , w3717 );
and ( w3719 , w3718 , w2582 );
not ( w3720 , w3719 );
and ( w3721 , w3720 , w2587 );
nor ( w3722 , w3721 , w2575 );
and ( w3723 , w3722 , w6110 );
not ( w3724 , w3620 );
and ( w3725 , w3724 , w3723 );
nor ( w3726 , w3725 , w312 );
and ( w3727 , w3726 , w12498 );
nor ( w3728 , w39 , w2674 );
and ( w3729 , w3728 , w5370 );
nor ( w3730 , w3729 , w43 );
nor ( w3731 , w3730 , w2735 );
and ( w3732 , w3731 , w2587 );
nor ( w3733 , w3732 , w2575 );
and ( w3734 , w3733 , w6110 );
nor ( w3735 , w3734 , w3113 );
nor ( w3736 , w3735 , w20 );
and ( w3737 , w3736 , w12142 );
and ( w3738 , w3737 , w8640 );
and ( w3739 , w3738 , w3106 );
and ( w3740 , w12921 , w3739 );
nor ( w3741 , w3740 , w2735 );
and ( w3742 , w3741 , w2624 );
and ( w3743 , w3742 , w2587 );
nor ( w3744 , w3743 , w2575 );
and ( w3745 , w12717 , w3744 );
and ( w3746 , w255 , w8848 );
not ( w3747 , w3746 );
and ( w3748 , w3747 , w3615 );
nor ( w3749 , w3748 , w384 );
and ( w3750 , w3749 , w12037 );
and ( w3751 , w3750 , w11166 );
and ( w3752 , w3751 , w5968 );
not ( w3753 , w3752 );
and ( w3754 , w3753 , w2582 );
not ( w3755 , w3754 );
and ( w3756 , w3755 , w2587 );
nor ( w3757 , w3756 , w2575 );
nor ( w3758 , w3745 , w3757 );
nor ( w3759 , w3758 , w310 );
nor ( w3760 , w3759 , w384 );
and ( w3761 , w3760 , w12037 );
nor ( w3762 , w2666 , w45 );
not ( w3763 , w3762 );
and ( w3764 , w3763 , w2664 );
nor ( w3765 , w35 , w2664 );
not ( w3766 , w3765 );
and ( w3767 , w3766 , w2666 );
nor ( w3768 , w3767 , w45 );
and ( w3769 , w3768 , w2587 );
not ( w3770 , w3769 );
and ( w3771 , w3770 , w2664 );
and ( w3772 , w3764 , w3771 );
and ( w3773 , w3772 , w2976 );
and ( w3774 , w3773 , w11166 );
nor ( w3775 , w3774 , w18 );
and ( w3776 , w3775 , w11166 );
and ( w3777 , w12921 , w3776 );
and ( w3778 , w3777 , w2587 );
not ( w3779 , w3778 );
and ( w3780 , w3779 , w2664 );
nor ( w3781 , w20 , w3780 );
and ( w3782 , w3781 , w2587 );
not ( w3783 , w3782 );
and ( w3784 , w3783 , w2664 );
and ( w3785 , w3734 , w3784 );
and ( w3786 , w3785 , w12142 );
nor ( w3787 , w3786 , w3116 );
nor ( w3788 , w3787 , w377 );
nor ( w3789 , w3788 , w3696 );
not ( w3790 , w3789 );
and ( w3791 , w3790 , w3417 );
nor ( w3792 , w3791 , w377 );
and ( w3793 , w3324 , w3833 );
nor ( w3794 , w3793 , w48 );
nor ( w3795 , w3794 , w105 );
and ( w3796 , w3795 , w12919 );
nor ( w3797 , w2615 , g10 );
not ( w3798 , w3796 );
and ( w3799 , w3798 , w3797 );
and ( w3800 , w3799 , w13477 );
and ( w3801 , w2664 , w45 );
and ( w3802 , w2664 , w6110 );
not ( w3803 , w239 );
and ( w3804 , w3802 , w3803 );
and ( w3805 , w3804 , w12424 );
nor ( w3806 , w3805 , w39 );
not ( w3807 , w3806 );
and ( w3808 , w3807 , w3802 );
and ( w3809 , w11140 , w2604 );
and ( w3810 , w3809 , w3802 );
not ( w3811 , w274 );
and ( w3812 , w3810 , w3811 );
and ( w3813 , w3812 , w8363 );
and ( w3814 , w3813 , w7485 );
and ( w3815 , w3814 , w12424 );
and ( w3816 , w3815 , w12144 );
not ( w3817 , w3816 );
and ( w3818 , w3817 , w2624 );
not ( w3819 , w3818 );
and ( w3820 , w3819 , w2573 );
and ( w3821 , w3820 , w6110 );
nor ( w3822 , w3808 , w3821 );
nor ( w3823 , w3822 , w41 );
and ( w3824 , w3823 , w12144 );
and ( w3825 , w3824 , w2573 );
and ( w3826 , w3825 , w6110 );
nor ( w3827 , w3801 , w3826 );
nor ( w3828 , w3827 , w43 );
not ( w3829 , w3324 );
and ( w3830 , w3828 , w3829 );
and ( w3831 , w3830 , w2976 );
nor ( w3832 , w3831 , w18 );
not ( w3833 , w3231 );
and ( w3834 , w3832 , w3833 );
nor ( w3835 , w3834 , w48 );
nor ( w3836 , w105 , w3835 );
not ( w3837 , w3836 );
and ( w3838 , w3837 , w19 );
and ( w3839 , w3838 , g11 );
and ( w3840 , w3839 , w2573 );
and ( w3841 , w3840 , w6110 );
nor ( w3842 , w3800 , w3841 );
and ( w3843 , w12921 , w3842 );
not ( w3844 , w3843 );
and ( w3845 , w3844 , w2573 );
and ( w3846 , w3845 , w6110 );
and ( w3847 , w12142 , w3846 );
nor ( w3848 , w3847 , w105 );
and ( w3849 , w3848 , w485 );
nor ( w3850 , w3849 , w2618 );
nor ( w3851 , w3850 , w18 );
and ( w3852 , w3851 , w8848 );
not ( w3853 , w3852 );
and ( w3854 , w3853 , w2582 );
not ( w3855 , w3854 );
and ( w3856 , w3855 , w2624 );
not ( w3857 , w3856 );
and ( w3858 , w3857 , w2573 );
and ( w3859 , w3858 , w6110 );
and ( w3860 , w3098 , w3859 );
not ( w3861 , w3860 );
and ( w3862 , w384 , w3861 );
not ( w3863 , w3862 );
and ( w3864 , w3863 , w2582 );
and ( w3865 , w3864 , w2573 );
and ( w3866 , w3865 , w6110 );
and ( w3867 , w12080 , w377 );
not ( w3868 , w3866 );
and ( w3869 , w3868 , w3867 );
and ( w3870 , w3869 , w377 );
not ( w3871 , w3870 );
and ( w3872 , w3871 , w2582 );
not ( w3873 , w3872 );
and ( w3874 , w3873 , w2587 );
nor ( w3875 , w3874 , w2575 );
not ( w3876 , w3792 );
and ( w3877 , w3876 , w3875 );
nor ( w3878 , w20 , w3877 );
nor ( w3879 , w3878 , w19 );
not ( w3880 , w3879 );
and ( w3881 , w3880 , g33 );
and ( w3882 , w3881 , w5968 );
not ( w3883 , w3882 );
and ( w3884 , w3883 , w2582 );
not ( w3885 , w3884 );
and ( w3886 , w3885 , w2624 );
and ( w3887 , w3886 , w2587 );
nor ( w3888 , w3887 , w2575 );
and ( w3889 , w3888 , w6110 );
and ( w3890 , w12921 , w3889 );
nor ( w3891 , w3890 , w3522 );
nor ( w3892 , w45 , w105 );
and ( w3893 , w3892 , w13477 );
and ( w3894 , w3893 , w11261 );
and ( w3895 , w3894 , w13477 );
nor ( w3896 , w45 , w2616 );
and ( w3897 , w3896 , w11166 );
nor ( w3898 , w3895 , w3897 );
nor ( w3899 , w3898 , w18 );
not ( w3900 , w2610 );
and ( w3901 , w3900 , w3899 );
nor ( w3902 , w3901 , w48 );
and ( w3903 , w3902 , w12144 );
nor ( w3904 , w3903 , w105 );
and ( w3905 , w3904 , w13477 );
and ( w3906 , w3905 , w11261 );
and ( w3907 , w3906 , w13477 );
and ( w3908 , w2605 , w3899 );
nor ( w3909 , w3908 , w41 );
not ( w3910 , w3909 );
and ( w3911 , w3910 , w3899 );
nor ( w3912 , w3911 , w48 );
nor ( w3913 , w3912 , w2616 );
nor ( w3914 , w3913 , w43 );
nor ( w3915 , w3914 , w2616 );
and ( w3916 , w3915 , w11166 );
and ( w3917 , w3916 , w12919 );
nor ( w3918 , w3907 , w3917 );
nor ( w3919 , w3918 , w18 );
and ( w3920 , w2615 , w11797 );
and ( w3921 , w3920 , w11533 );
nor ( w3922 , w3921 , g12 );
and ( w3923 , w3922 , w11797 );
nor ( w3924 , w3923 , w105 );
and ( w3925 , w3924 , w20 );
nor ( w3926 , w3919 , w3925 );
not ( w3927 , w3926 );
and ( w3928 , w3927 , g29 );
and ( w3929 , w3928 , g28 );
not ( w3930 , w3929 );
and ( w3931 , w3930 , g28 );
not ( w3932 , w3931 );
and ( w3933 , w3932 , g29 );
not ( w3934 , w3933 );
and ( w3935 , w3934 , g29 );
nor ( w3936 , w3935 , w134 );
and ( w3937 , w3936 , w2908 );
and ( w3938 , w3937 , g29 );
not ( w3939 , w3938 );
and ( w3940 , w3939 , w3417 );
nor ( w3941 , w3940 , w19 );
not ( w3942 , w3941 );
and ( w3943 , w3942 , w20 );
and ( w3944 , w3943 , w11166 );
not ( w3945 , w3944 );
and ( w3946 , w3945 , w20 );
not ( w3947 , w2961 );
and ( w3948 , w3946 , w3947 );
nor ( w3949 , w134 , g28 );
nor ( w3950 , w3949 , g28 );
not ( w3951 , w3950 );
and ( w3952 , w3951 , g29 );
and ( w3953 , w2908 , g28 );
not ( w3954 , w3953 );
and ( w3955 , w3954 , g28 );
nor ( w3956 , w3955 , g29 );
nor ( w3957 , w3952 , w3956 );
nor ( w3958 , w3957 , w255 );
not ( w3959 , w3958 );
and ( w3960 , w3959 , w3097 );
and ( w3961 , w3960 , w8640 );
and ( w3962 , w3961 , w19 );
nor ( w3963 , w3962 , w3417 );
and ( w3964 , w3937 , w13206 );
and ( w3965 , w3964 , w12199 );
and ( w3966 , w3965 , w13206 );
and ( w3967 , w3966 , w12717 );
and ( w3968 , w3952 , w12080 );
and ( w3969 , w3968 , g29 );
nor ( w3970 , w3967 , w3969 );
not ( w3971 , w3970 );
and ( w3972 , w3971 , g29 );
nor ( w3973 , w3972 , w3956 );
nor ( w3974 , w3973 , w377 );
and ( w3975 , w3974 , w2587 );
not ( w3976 , w3975 );
and ( w3977 , w3976 , w2664 );
and ( w3978 , w3977 , w3784 );
and ( w3979 , w3978 , w6110 );
not ( w3980 , w3963 );
and ( w3981 , w3980 , w3979 );
and ( w3982 , w3981 , w12921 );
and ( w3983 , w3982 , w2976 );
nor ( w3984 , w3983 , w20 );
and ( w3985 , w3984 , w5597 );
nor ( w3986 , w3985 , w105 );
and ( w3987 , w3986 , w12498 );
nor ( w3988 , w3987 , w2961 );
and ( w3989 , w3988 , w12498 );
and ( w3990 , w3989 , g33 );
and ( w3991 , w12717 , w3990 );
not ( w3992 , w3991 );
and ( w3993 , w3992 , w2582 );
not ( w3994 , w3993 );
and ( w3995 , w3994 , w2624 );
not ( w3996 , w3995 );
and ( w3997 , w3996 , w2573 );
and ( w3998 , w3997 , w6110 );
not ( w3999 , w3948 );
and ( w4000 , w3999 , w3998 );
not ( w4001 , w3867 );
and ( w4002 , w4000 , w4001 );
and ( w4003 , w20 , w3924 );
not ( w4004 , w4003 );
and ( w4005 , w4004 , w3866 );
not ( w4006 , w4005 );
and ( w4007 , w377 , w4006 );
and ( w4008 , w255 , w3925 );
not ( w4009 , w4008 );
and ( w4010 , w4009 , w3417 );
nor ( w4011 , w4010 , w19 );
and ( w4012 , w20 , w4011 );
not ( w4013 , w4012 );
and ( w4014 , w4013 , w3998 );
nor ( w4015 , w377 , w4014 );
and ( w4016 , w4015 , w384 );
and ( w4017 , w4016 , g33 );
and ( w4018 , w4017 , w12717 );
not ( w4019 , w4018 );
and ( w4020 , w4019 , w2582 );
not ( w4021 , w4020 );
and ( w4022 , w4021 , w2624 );
not ( w4023 , w4022 );
and ( w4024 , w4023 , w2573 );
and ( w4025 , w4024 , w6110 );
not ( w4026 , w4007 );
and ( w4027 , w4026 , w4025 );
not ( w4028 , w4027 );
and ( w4029 , w384 , w4028 );
and ( w4030 , w4029 , g33 );
and ( w4031 , w12717 , w4030 );
not ( w4032 , w4031 );
and ( w4033 , w4032 , w2582 );
not ( w4034 , w4033 );
and ( w4035 , w4034 , w2624 );
not ( w4036 , w4035 );
and ( w4037 , w4036 , w2573 );
and ( w4038 , w4037 , w6110 );
nor ( w4039 , w4002 , w4038 );
and ( w4040 , w4039 , w384 );
and ( w4041 , w3925 , w377 );
and ( w4042 , w4041 , w12080 );
and ( w4043 , w4042 , w12717 );
not ( w4044 , w4043 );
and ( w4045 , w4044 , w2582 );
not ( w4046 , w4045 );
and ( w4047 , w4046 , w2624 );
not ( w4048 , w4047 );
and ( w4049 , w4048 , w3417 );
nor ( w4050 , w4049 , w19 );
not ( w4051 , w4050 );
and ( w4052 , w4051 , w3427 );
not ( w4053 , w4052 );
and ( w4054 , w20 , w4053 );
not ( w4055 , w2618 );
and ( w4056 , w4055 , w2976 );
and ( w4057 , w4056 , w3097 );
nor ( w4058 , w4057 , w3113 );
and ( w4059 , w12921 , w4058 );
not ( w4060 , w4059 );
and ( w4061 , w4060 , w2582 );
not ( w4062 , w4061 );
and ( w4063 , w4062 , w2624 );
not ( w4064 , w4063 );
and ( w4065 , w4064 , w2573 );
and ( w4066 , w4065 , w6110 );
not ( w4067 , w3849 );
and ( w4068 , w4067 , w4066 );
not ( w4069 , w4068 );
and ( w4070 , w4069 , w377 );
not ( w4071 , w4070 );
and ( w4072 , w4071 , w3417 );
and ( w4073 , w4072 , w8848 );
and ( w4074 , w4073 , w12921 );
nor ( w4075 , w4074 , w19 );
and ( w4076 , w4075 , w12921 );
and ( w4077 , w3780 , w2922 );
nor ( w4078 , w20 , w4077 );
not ( w4079 , w4078 );
and ( w4080 , w4079 , w2582 );
not ( w4081 , w4080 );
and ( w4082 , w4081 , w2624 );
not ( w4083 , w4082 );
and ( w4084 , w4083 , w2573 );
and ( w4085 , w4084 , w6110 );
nor ( w4086 , w105 , w4085 );
not ( w4087 , w4086 );
and ( w4088 , w4087 , w2976 );
and ( w4089 , w4088 , w12921 );
and ( w4090 , w4089 , w3097 );
nor ( w4091 , w4090 , w3113 );
and ( w4092 , w4091 , w12921 );
and ( w4093 , w12717 , w4092 );
and ( w4094 , w4093 , w2624 );
not ( w4095 , w4094 );
and ( w4096 , w4095 , w2573 );
and ( w4097 , w4096 , w6110 );
nor ( w4098 , w310 , w4097 );
not ( w4099 , w4098 );
and ( w4100 , w4099 , w2573 );
and ( w4101 , w4100 , w6110 );
nor ( w4102 , w35 , w4101 );
not ( w4103 , w4102 );
and ( w4104 , w4103 , w2666 );
nor ( w4105 , w4104 , w45 );
nor ( w4106 , w4105 , w20 );
and ( w4107 , w4106 , w3097 );
nor ( w4108 , w4107 , w20 );
and ( w4109 , w12717 , w4108 );
not ( w4110 , w4109 );
and ( w4111 , w4110 , w2582 );
not ( w4112 , w4111 );
and ( w4113 , w4112 , w2624 );
not ( w4114 , w4113 );
and ( w4115 , w4114 , w2573 );
and ( w4116 , w4115 , w6110 );
and ( w4117 , w4116 , w2688 );
nor ( w4118 , w105 , w4117 );
not ( w4119 , w4118 );
and ( w4120 , w4119 , w2976 );
and ( w4121 , w4120 , w12921 );
and ( w4122 , w4121 , w3097 );
nor ( w4123 , w4122 , w3113 );
and ( w4124 , w4123 , w12921 );
and ( w4125 , w12717 , w4124 );
not ( w4126 , w4125 );
and ( w4127 , w4126 , w2582 );
not ( w4128 , w4127 );
and ( w4129 , w4128 , w2624 );
not ( w4130 , w4129 );
and ( w4131 , w4130 , w2573 );
and ( w4132 , w4131 , w3427 );
nor ( w4133 , w310 , w4132 );
not ( w4134 , w4133 );
and ( w4135 , w4134 , w2582 );
and ( w4136 , w4135 , w2573 );
and ( w4137 , w4136 , w6110 );
not ( w4138 , w4076 );
and ( w4139 , w4138 , w4137 );
nor ( w4140 , w4139 , w255 );
and ( w4141 , w4140 , g33 );
and ( w4142 , w12717 , w4141 );
not ( w4143 , w4142 );
and ( w4144 , w4143 , w2582 );
not ( w4145 , w4144 );
and ( w4146 , w4145 , w2624 );
not ( w4147 , w4146 );
and ( w4148 , w4147 , w2573 );
not ( w4149 , w4054 );
and ( w4150 , w4149 , w4148 );
and ( w4151 , w2573 , w105 );
and ( w4152 , w4151 , w2961 );
not ( w4153 , w4152 );
and ( w4154 , w105 , w4153 );
and ( w4155 , w12717 , w4154 );
not ( w4156 , w4155 );
and ( w4157 , w4156 , w2582 );
not ( w4158 , w4157 );
and ( w4159 , w4158 , w2624 );
not ( w4160 , w4159 );
and ( w4161 , w4160 , w2573 );
and ( w4162 , w4161 , w6110 );
and ( w4163 , w4150 , w4162 );
nor ( w4164 , w4163 , w255 );
and ( w4165 , w4164 , g33 );
and ( w4166 , w12717 , w4165 );
not ( w4167 , w4166 );
and ( w4168 , w4167 , w2582 );
and ( w4169 , w4168 , w2573 );
and ( w4170 , w4169 , w6110 );
not ( w4171 , w4040 );
and ( w4172 , w4171 , w4170 );
not ( w4173 , w4172 );
and ( w4174 , w4173 , g33 );
not ( w4175 , w4174 );
and ( w4176 , w4175 , w3582 );
not ( w4177 , w4176 );
and ( w4178 , w4177 , g32 );
and ( w4179 , w3 , g5 );
nor ( w4180 , w4179 , w2553 );
not ( w4181 , w4180 );
and ( w4182 , w4181 , g47 );
nor ( w4183 , w4182 , w2647 );
nor ( w4184 , w4178 , w4183 );
nor ( w4185 , w4184 , w310 );
not ( w4186 , w3577 );
and ( w4187 , w4185 , w4186 );
not ( w4188 , w4187 );
and ( w4189 , w4188 , w2582 );
not ( w4190 , w4189 );
and ( w4191 , w4190 , w2624 );
not ( w4192 , w4191 );
and ( w4193 , w4192 , w2573 );
and ( w4194 , w4193 , w6110 );
not ( w4195 , w4194 );
and ( w4196 , w4195 , g33 );
nor ( w4197 , w3891 , w4196 );
nor ( w4198 , w310 , w3431 );
not ( w4199 , w4198 );
and ( w4200 , w4199 , w2587 );
and ( w4201 , w4197 , w5649 );
and ( w4202 , w4201 , w384 );
and ( w4203 , w12142 , w2680 );
not ( w4204 , w4203 );
and ( w4205 , w4204 , w2624 );
not ( w4206 , w2628 );
and ( w4207 , w4206 , w4205 );
and ( w4208 , w4207 , w12919 );
and ( w4209 , w4208 , w11166 );
and ( w4210 , w2573 , w2664 );
nor ( w4211 , w20 , w4210 );
not ( w4212 , w4211 );
and ( w4213 , w4212 , w2582 );
not ( w4214 , w4213 );
and ( w4215 , w4214 , w2624 );
not ( w4216 , w4215 );
and ( w4217 , w4216 , w2573 );
and ( w4218 , w4217 , w6110 );
not ( w4219 , w4209 );
and ( w4220 , w4219 , w4218 );
not ( w4221 , w4220 );
and ( w4222 , w4221 , w485 );
nor ( w4223 , w4222 , w20 );
and ( w4224 , w4223 , w4066 );
nor ( w4225 , w4224 , w20 );
not ( w4226 , w4225 );
and ( w4227 , w4226 , w2582 );
not ( w4228 , w4227 );
and ( w4229 , w4228 , w2624 );
and ( w4230 , w4229 , w2587 );
nor ( w4231 , w4230 , w2575 );
and ( w4232 , w4231 , w6110 );
and ( w4233 , w12921 , w4232 );
and ( w4234 , w4218 , w12921 );
and ( w4235 , w4234 , w105 );
not ( w4236 , w4235 );
and ( w4237 , w4236 , g13 );
not ( w4238 , w4237 );
and ( w4239 , w4238 , g13 );
nor ( w4240 , w4239 , w2735 );
and ( w4241 , w4240 , w2624 );
and ( w4242 , w4241 , w2587 );
nor ( w4243 , w4242 , w2575 );
nor ( w4244 , w4233 , w4243 );
not ( w4245 , w4170 );
and ( w4246 , w4245 , w2587 );
nor ( w4247 , w4246 , w2575 );
not ( w4248 , w4244 );
and ( w4249 , w4248 , w4247 );
nor ( w4250 , w4249 , g29 );
and ( w4251 , w4250 , w3867 );
and ( w4252 , w4251 , w377 );
not ( w4253 , w4252 );
and ( w4254 , w4253 , w3696 );
and ( w4255 , w8640 , w4066 );
and ( w4256 , w4255 , w12921 );
nor ( w4257 , w4256 , w4243 );
not ( w4258 , w4257 );
and ( w4259 , w4258 , w4247 );
nor ( w4260 , w4259 , g29 );
and ( w4261 , w4260 , w3867 );
and ( w4262 , w4261 , w377 );
nor ( w4263 , w3734 , w3116 );
nor ( w4264 , w20 , w4263 );
and ( w4265 , w4264 , w6110 );
and ( w4266 , w4265 , w12142 );
and ( w4267 , w4266 , w11166 );
and ( w4268 , w4267 , w12498 );
and ( w4269 , w4268 , w3417 );
nor ( w4270 , w4269 , w2961 );
and ( w4271 , w4270 , w12498 );
and ( w4272 , w4271 , w5968 );
and ( w4273 , w4272 , w2624 );
and ( w4274 , w4273 , w2587 );
nor ( w4275 , w4274 , w2575 );
and ( w4276 , w4275 , w6110 );
not ( w4277 , w4262 );
and ( w4278 , w4277 , w4276 );
and ( w4279 , w4278 , w8848 );
nor ( w4280 , w4279 , w310 );
and ( w4281 , w4280 , g33 );
and ( w4282 , w4281 , w5968 );
not ( w4283 , w4282 );
and ( w4284 , w4283 , w2582 );
not ( w4285 , w4284 );
and ( w4286 , w4285 , w2587 );
nor ( w4287 , w4286 , w2575 );
and ( w4288 , w4287 , w6110 );
nor ( w4289 , w4254 , w4288 );
and ( w4290 , w8848 , w4289 );
not ( w4291 , w4290 );
and ( w4292 , w4291 , w3506 );
and ( w4293 , w4292 , w11852 );
nor ( w4294 , w4293 , w310 );
and ( w4295 , w4294 , g33 );
and ( w4296 , w4295 , w5968 );
not ( w4297 , w4296 );
and ( w4298 , w4297 , w2582 );
not ( w4299 , w4298 );
and ( w4300 , w4299 , w2587 );
nor ( w4301 , w4300 , w2575 );
and ( w4302 , w4301 , w6110 );
nor ( w4303 , w4202 , w4302 );
and ( w4304 , w4303 , w12717 );
not ( w4305 , w3597 );
and ( w4306 , w4304 , w4305 );
not ( w4307 , w4306 );
and ( w4308 , w4307 , w3582 );
not ( w4309 , w4308 );
and ( w4310 , w4309 , g33 );
not ( w4311 , w4310 );
and ( w4312 , w4311 , w2647 );
not ( w4313 , w4312 );
and ( w4314 , w4313 , g32 );
not ( w4315 , w4314 );
and ( w4316 , w4315 , g32 );
and ( w4317 , w4316 , g33 );
nor ( w4318 , w4317 , w2735 );
not ( w4319 , w4318 );
and ( w4320 , w4319 , w2582 );
not ( w4321 , w4320 );
and ( w4322 , w4321 , w2624 );
and ( w4323 , w4322 , w2587 );
nor ( w4324 , w4323 , w2575 );
and ( w4325 , w4324 , w6110 );
and ( w4326 , w4325 , w2758 );
and ( w4327 , w4326 , w2573 );
and ( w4328 , w4327 , w2664 );
and ( w4329 , w4328 , w12921 );
and ( w4330 , w4329 , w3734 );
and ( w4331 , w4330 , w12142 );
and ( w4332 , w12921 , w4331 );
nor ( w4333 , w2605 , w41 );
not ( w4334 , w4333 );
and ( w4335 , w4334 , w3222 );
and ( w4336 , w3163 , w2605 );
and ( w4337 , w4336 , w11347 );
and ( w4338 , w4337 , w239 );
nor ( w4339 , w2672 , w4338 );
nor ( w4340 , w4339 , w255 );
nor ( w4341 , w4340 , w41 );
not ( w4342 , w4341 );
and ( w4343 , w4335 , w4342 );
and ( w4344 , w4343 , w8848 );
nor ( w4345 , w4344 , w3958 );
nor ( w4346 , w4345 , g31 );
and ( w4347 , w4346 , w12199 );
and ( w4348 , w4347 , w13206 );
and ( w4349 , w4348 , w3324 );
nor ( w4350 , w377 , w3297 );
nor ( w4351 , w4350 , w105 );
nor ( w4352 , w20 , w4351 );
and ( w4353 , w12717 , w4352 );
nor ( w4354 , w4349 , w4353 );
and ( w4355 , w8363 , w2592 );
not ( w4356 , w4355 );
and ( w4357 , w4356 , w2664 );
nor ( w4358 , w20 , w4357 );
not ( w4359 , w4358 );
and ( w4360 , w4359 , w2573 );
and ( w4361 , w4360 , w6110 );
and ( w4362 , w4354 , w4361 );
nor ( w4363 , w4362 , w39 );
not ( w4364 , w4363 );
and ( w4365 , w4364 , w2666 );
nor ( w4366 , w4365 , w45 );
not ( w4367 , w4366 );
and ( w4368 , w4367 , w2664 );
nor ( w4369 , w4368 , w48 );
and ( w4370 , w11166 , w4369 );
not ( w4371 , w4370 );
and ( w4372 , w4371 , w2976 );
and ( w4373 , w4372 , w2573 );
nor ( w4374 , w4373 , w3113 );
and ( w4375 , w12921 , w4374 );
and ( w4376 , w12498 , w4375 );
and ( w4377 , w4376 , g33 );
and ( w4378 , w12717 , w4377 );
and ( w4379 , w4378 , w12080 );
and ( w4380 , w4379 , w2624 );
not ( w4381 , w4380 );
and ( w4382 , w4381 , w2573 );
and ( w4383 , w4382 , w6110 );
and ( w4384 , w4383 , w384 );
and ( w4385 , w4384 , w13206 );
and ( w4386 , w4385 , w8640 );
and ( w4387 , w4386 , w19 );
nor ( w4388 , w4387 , w3417 );
and ( w4389 , w4388 , w12498 );
and ( w4390 , w12717 , w4389 );
and ( w4391 , w4390 , w12080 );
not ( w4392 , w4391 );
and ( w4393 , w4392 , w2573 );
and ( w4394 , w4393 , w6110 );
and ( w4395 , w4394 , w3597 );
nor ( w4396 , w4395 , w3575 );
and ( w4397 , w4396 , g32 );
not ( w4398 , w4397 );
and ( w4399 , w4398 , g32 );
and ( w4400 , w4399 , w5094 );
and ( w4401 , w4400 , g33 );
and ( w4402 , w4401 , w312 );
nor ( w4403 , w4402 , w2735 );
not ( w4404 , w4403 );
and ( w4405 , w4404 , w2582 );
not ( w4406 , w4405 );
and ( w4407 , w4406 , w2624 );
and ( w4408 , w4407 , w2587 );
nor ( w4409 , w4408 , w2575 );
and ( w4410 , w4409 , w6110 );
nor ( w4411 , w377 , w4410 );
not ( w4412 , w4411 );
and ( w4413 , w4412 , w312 );
nor ( w4414 , w4413 , w2735 );
not ( w4415 , w4414 );
and ( w4416 , w4415 , w2582 );
not ( w4417 , w4416 );
and ( w4418 , w4417 , w2587 );
nor ( w4419 , w4418 , w2575 );
and ( w4420 , w4325 , w4419 );
and ( w4421 , w4420 , w3615 );
and ( w4422 , w4421 , w312 );
nor ( w4423 , w4422 , w2735 );
not ( w4424 , w4423 );
and ( w4425 , w4424 , w2582 );
not ( w4426 , w4425 );
and ( w4427 , w4426 , w2587 );
nor ( w4428 , w4427 , w2575 );
and ( w4429 , w4428 , w19 );
and ( w4430 , g31 , w11852 );
and ( w4431 , w4430 , w310 );
and ( w4432 , w3623 , w255 );
and ( w4433 , w4432 , w8848 );
not ( w4434 , w4433 );
and ( w4435 , w4434 , w3615 );
nor ( w4436 , w4435 , w3696 );
and ( w4437 , w4436 , w12498 );
not ( w4438 , w3744 );
and ( w4439 , w4437 , w4438 );
and ( w4440 , w4439 , w12717 );
and ( w4441 , w4440 , w11852 );
and ( w4442 , w4441 , w11166 );
and ( w4443 , w4442 , w5968 );
not ( w4444 , w4443 );
and ( w4445 , w4444 , w2582 );
not ( w4446 , w4445 );
and ( w4447 , w4446 , w2587 );
nor ( w4448 , w4447 , w2575 );
and ( w4449 , w4448 , w2582 );
not ( w4450 , w4449 );
and ( w4451 , w4450 , w2587 );
nor ( w4452 , w4451 , w2575 );
not ( w4453 , w4431 );
and ( w4454 , w4453 , w4452 );
nor ( w4455 , w4454 , w105 );
and ( w4456 , w4455 , w12532 );
and ( w4457 , w4456 , w5968 );
not ( w4458 , w4457 );
and ( w4459 , w4458 , w2582 );
not ( w4460 , w4459 );
and ( w4461 , w4460 , w2587 );
nor ( w4462 , w4461 , w2575 );
and ( w4463 , w12037 , w4462 );
not ( w4464 , w3486 );
and ( w4465 , w4464 , g32 );
not ( w4466 , w4465 );
and ( w4467 , w4466 , g32 );
and ( w4468 , w4467 , w5094 );
and ( w4469 , w4468 , g33 );
and ( w4470 , w4469 , w312 );
and ( w4471 , w4470 , w12717 );
nor ( w4472 , w4471 , w2994 );
and ( w4473 , w4472 , w11166 );
and ( w4474 , w4473 , w12532 );
and ( w4475 , w4474 , w5968 );
not ( w4476 , w4475 );
and ( w4477 , w4476 , w2582 );
not ( w4478 , w4477 );
and ( w4479 , w4478 , w2624 );
and ( w4480 , w4479 , w2587 );
nor ( w4481 , w4480 , w2575 );
nor ( w4482 , w4463 , w4481 );
nor ( w4483 , w4482 , w19 );
and ( w4484 , w4483 , w12080 );
nor ( w4485 , w4484 , w2735 );
not ( w4486 , w4485 );
and ( w4487 , w4486 , w2582 );
not ( w4488 , w4487 );
and ( w4489 , w4488 , w2587 );
nor ( w4490 , w4489 , w2575 );
nor ( w4491 , w4454 , w308 );
and ( w4492 , w4491 , w5968 );
not ( w4493 , w4492 );
and ( w4494 , w4493 , w2582 );
not ( w4495 , w4494 );
and ( w4496 , w4495 , w2587 );
nor ( w4497 , w4496 , w2575 );
and ( w4498 , w12037 , w4497 );
nor ( w4499 , w4498 , w2735 );
not ( w4500 , w4499 );
and ( w4501 , w4500 , w2582 );
not ( w4502 , w4501 );
and ( w4503 , w4502 , w2587 );
nor ( w4504 , w4503 , w2575 );
nor ( w4505 , w4490 , w4504 );
and ( w4506 , w4505 , w5898 );
and ( w4507 , w4506 , w11166 );
and ( w4508 , w4507 , w5968 );
not ( w4509 , w4508 );
and ( w4510 , w4509 , w2582 );
not ( w4511 , w4510 );
and ( w4512 , w4511 , w2587 );
nor ( w4513 , w4512 , w2575 );
nor ( w4514 , w4429 , w4513 );
nor ( w4515 , w4514 , w384 );
not ( w4516 , w4515 );
and ( w4517 , w4516 , g31 );
and ( w4518 , w4517 , w11852 );
and ( w4519 , w4518 , w310 );
not ( w4520 , w4519 );
and ( w4521 , w4520 , w3605 );
not ( w4522 , w4521 );
and ( w4523 , w4522 , g32 );
and ( w4524 , w4523 , g33 );
not ( w4525 , w2745 );
and ( w4526 , w4525 , w2752 );
and ( w4527 , w4526 , w2758 );
and ( w4528 , w4527 , w2573 );
and ( w4529 , w4528 , w2664 );
and ( w4530 , w4529 , w12921 );
and ( w4531 , w4530 , w3734 );
and ( w4532 , w4531 , w12142 );
and ( w4533 , w12921 , w4532 );
nor ( w4534 , w4533 , w4513 );
and ( w4535 , w4534 , w8848 );
and ( w4536 , w2589 , w3615 );
and ( w4537 , w4536 , w4452 );
nor ( w4538 , w4537 , w308 );
and ( w4539 , w4538 , w5968 );
not ( w4540 , w4539 );
and ( w4541 , w4540 , w2582 );
not ( w4542 , w4541 );
and ( w4543 , w4542 , w2587 );
nor ( w4544 , w4543 , w2575 );
and ( w4545 , w3615 , w4544 );
and ( w4546 , w4545 , w4452 );
nor ( w4547 , w4546 , w312 );
and ( w4548 , w4547 , w12532 );
and ( w4549 , w4548 , w5968 );
not ( w4550 , w4549 );
and ( w4551 , w4550 , w2582 );
not ( w4552 , w4551 );
and ( w4553 , w4552 , w2587 );
nor ( w4554 , w4553 , w2575 );
not ( w4555 , w4535 );
and ( w4556 , w4555 , w4554 );
not ( w4557 , w4556 );
and ( w4558 , w4557 , g31 );
and ( w4559 , w310 , w4558 );
not ( w4560 , w4559 );
and ( w4561 , w4560 , w4452 );
nor ( w4562 , w4561 , w312 );
and ( w4563 , w4562 , w11852 );
and ( w4564 , w4563 , w5898 );
and ( w4565 , w4564 , w11166 );
and ( w4566 , w4565 , w12532 );
and ( w4567 , w4566 , w5968 );
not ( w4568 , w4567 );
and ( w4569 , w4568 , w2582 );
not ( w4570 , w4569 );
and ( w4571 , w4570 , w2624 );
and ( w4572 , w4571 , w2587 );
nor ( w4573 , w4572 , w2575 );
and ( w4574 , w4573 , w6110 );
not ( w4575 , w4524 );
and ( w4576 , w4575 , w4574 );
nor ( w4577 , w4576 , w4504 );
and ( w4578 , w4577 , w12532 );
and ( w4579 , w4578 , w5968 );
not ( w4580 , w4579 );
and ( w4581 , w4580 , w2582 );
not ( w4582 , w4581 );
and ( w4583 , w4582 , w2587 );
nor ( w4584 , w4583 , w2575 );
nor ( w4585 , w4332 , w4584 );
and ( w4586 , w4585 , g32 );
and ( w4587 , w4586 , g33 );
not ( w4588 , w4587 );
and ( w4589 , w4588 , w4574 );
nor ( w4590 , w4589 , w4504 );
and ( w4591 , w4590 , w5898 );
and ( w4592 , w4591 , w11166 );
and ( w4593 , w4592 , w5968 );
not ( w4594 , w4593 );
and ( w4595 , w4594 , w2582 );
not ( w4596 , w4595 );
and ( w4597 , w4596 , w2624 );
and ( w4598 , w4597 , w2587 );
nor ( w4599 , w4598 , w2575 );
and ( w4600 , w4599 , w6110 );
not ( w4601 , w4600 );
and ( w4602 , w3761 , w4601 );
and ( w4603 , w4602 , w12532 );
and ( w4604 , w4603 , w5968 );
not ( w4605 , w4604 );
and ( w4606 , w4605 , w2582 );
not ( w4607 , w4606 );
and ( w4608 , w4607 , w2587 );
nor ( w4609 , w4608 , w2575 );
and ( w4610 , w12037 , w4609 );
nor ( w4611 , w4610 , w4600 );
and ( w4612 , w4611 , w5968 );
not ( w4613 , w4612 );
and ( w4614 , w4613 , w2582 );
not ( w4615 , w4614 );
and ( w4616 , w4615 , w2587 );
nor ( w4617 , w4616 , w2575 );
and ( w4618 , w3727 , w4950 );
and ( w4619 , w4618 , w5898 );
and ( w4620 , w4619 , w11166 );
and ( w4621 , w4620 , w12532 );
and ( w4622 , w4621 , w5968 );
not ( w4623 , w4622 );
and ( w4624 , w4623 , w2582 );
not ( w4625 , w4624 );
and ( w4626 , w4625 , w2587 );
nor ( w4627 , w4626 , w2575 );
and ( w4628 , w3611 , w4627 );
nor ( w4629 , w4628 , w2994 );
and ( w4630 , w4629 , w11166 );
and ( w4631 , w4630 , w5968 );
not ( w4632 , w4631 );
and ( w4633 , w4632 , w2582 );
not ( w4634 , w4633 );
and ( w4635 , w4634 , w2624 );
and ( w4636 , w4635 , w2587 );
nor ( w4637 , w4636 , w2575 );
not ( w4638 , w3157 );
and ( w4639 , w4638 , w4637 );
not ( w4640 , w4639 );
and ( w4641 , w4640 , g31 );
and ( w4642 , w4641 , w11852 );
and ( w4643 , w4642 , w310 );
not ( w4644 , w4643 );
and ( w4645 , w4644 , w3605 );
not ( w4646 , w4645 );
and ( w4647 , w4646 , w312 );
not ( w4648 , w4647 );
and ( w4649 , w4648 , w3615 );
and ( w4650 , w3151 , w310 );
not ( w4651 , w4650 );
and ( w4652 , w4651 , w3615 );
not ( w4653 , w4652 );
and ( w4654 , w4653 , w310 );
and ( w4655 , w4654 , w377 );
and ( w4656 , w4655 , w12080 );
and ( w4657 , w4656 , w11852 );
and ( w4658 , w377 , w4657 );
and ( w4659 , w4658 , w12037 );
and ( w4660 , w12717 , w3757 );
nor ( w4661 , w4660 , w4627 );
and ( w4662 , w4661 , w11852 );
and ( w4663 , w4662 , w12037 );
and ( w4664 , w4663 , w5898 );
and ( w4665 , w4664 , w11166 );
and ( w4666 , w4665 , w12532 );
and ( w4667 , w4666 , w5968 );
not ( w4668 , w4667 );
and ( w4669 , w4668 , w2582 );
not ( w4670 , w4669 );
and ( w4671 , w4670 , w2587 );
nor ( w4672 , w4671 , w2575 );
not ( w4673 , w4659 );
and ( w4674 , w4673 , w4672 );
not ( w4675 , w4674 );
and ( w4676 , w20 , w4675 );
and ( w4677 , w3431 , w2587 );
and ( w4678 , w4677 , w12080 );
not ( w4679 , w4678 );
and ( w4680 , w4679 , w2664 );
and ( w4681 , w4680 , w3683 );
and ( w4682 , w4681 , w2888 );
nor ( w4683 , w4682 , w3486 );
and ( w4684 , w4683 , g32 );
not ( w4685 , w4684 );
and ( w4686 , w4685 , g32 );
and ( w4687 , w4686 , g33 );
and ( w4688 , w4687 , w5094 );
not ( w4689 , w4688 );
and ( w4690 , w4689 , w312 );
and ( w4691 , w2890 , w2888 );
not ( w4692 , w4691 );
and ( w4693 , w4692 , w377 );
and ( w4694 , w4693 , w12080 );
and ( w4695 , w377 , w4694 );
and ( w4696 , w3643 , w12424 );
and ( w4697 , w4696 , w7803 );
nor ( w4698 , w4697 , w39 );
and ( w4699 , w4698 , w5370 );
nor ( w4700 , w4699 , w43 );
nor ( w4701 , w4700 , w2735 );
and ( w4702 , w4701 , w2587 );
nor ( w4703 , w4702 , w2575 );
and ( w4704 , w4703 , w6110 );
not ( w4705 , w4704 );
and ( w4706 , w4705 , w2587 );
nor ( w4707 , w4706 , w2575 );
and ( w4708 , w4707 , w6110 );
and ( w4709 , w3639 , w7803 );
nor ( w4710 , w4709 , w2680 );
and ( w4711 , w4710 , w11140 );
and ( w4712 , w4711 , w12117 );
nor ( w4713 , w4712 , w43 );
nor ( w4714 , w4713 , w2735 );
and ( w4715 , w4714 , w2587 );
nor ( w4716 , w4715 , w2575 );
and ( w4717 , w4716 , w6110 );
and ( w4718 , w4708 , w4717 );
and ( w4719 , w4718 , w8640 );
nor ( w4720 , w4719 , w3683 );
nor ( w4721 , w4720 , w2592 );
and ( w4722 , w4721 , w12921 );
and ( w4723 , w4722 , w12144 );
and ( w4724 , w4723 , w12142 );
and ( w4725 , w12921 , w4724 );
nor ( w4726 , w4725 , w19 );
nor ( w4727 , w4726 , w105 );
and ( w4728 , w4727 , w3615 );
nor ( w4729 , w4728 , w2961 );
and ( w4730 , w4729 , w12498 );
and ( w4731 , w4730 , w5898 );
and ( w4732 , w4731 , w11166 );
and ( w4733 , w4732 , w5968 );
not ( w4734 , w4733 );
and ( w4735 , w4734 , w2582 );
not ( w4736 , w4735 );
and ( w4737 , w4736 , w2624 );
and ( w4738 , w4737 , w2587 );
nor ( w4739 , w4738 , w2575 );
and ( w4740 , w4739 , w6110 );
not ( w4741 , w4695 );
and ( w4742 , w4741 , w4740 );
and ( w4743 , w4742 , w6110 );
not ( w4744 , w4743 );
and ( w4745 , w4744 , g31 );
and ( w4746 , w310 , w4745 );
nor ( w4747 , w3723 , w4617 );
and ( w4748 , w4747 , w12532 );
and ( w4749 , w4748 , w5968 );
not ( w4750 , w4749 );
and ( w4751 , w4750 , w2582 );
not ( w4752 , w4751 );
and ( w4753 , w4752 , w2587 );
nor ( w4754 , w4753 , w2575 );
not ( w4755 , w4746 );
and ( w4756 , w4755 , w4754 );
nor ( w4757 , w4756 , w384 );
and ( w4758 , w4757 , w12037 );
and ( w4759 , w4758 , w8848 );
and ( w4760 , w4759 , w485 );
nor ( w4761 , w3757 , w4754 );
nor ( w4762 , w4761 , w312 );
nor ( w4763 , w4762 , w3605 );
and ( w4764 , w4763 , w5048 );
not ( w4765 , w4764 );
and ( w4766 , w4765 , w3097 );
nor ( w4767 , w2778 , w2855 );
nor ( w4768 , w4767 , w35 );
and ( w4769 , w4768 , w7485 );
and ( w4770 , w4769 , w12424 );
and ( w4771 , w4770 , w7803 );
nor ( w4772 , w4771 , w39 );
and ( w4773 , w4772 , w5422 );
and ( w4774 , w4773 , w5370 );
nor ( w4775 , w4774 , w2592 );
and ( w4776 , w4775 , w12144 );
and ( w4777 , w4776 , w12142 );
nor ( w4778 , w20 , w4777 );
and ( w4779 , w4778 , w5968 );
not ( w4780 , w4779 );
and ( w4781 , w4780 , w2582 );
not ( w4782 , w4781 );
and ( w4783 , w4782 , w2624 );
and ( w4784 , w4783 , w2587 );
nor ( w4785 , w4784 , w2575 );
and ( w4786 , w4785 , w6110 );
not ( w4787 , w4786 );
and ( w4788 , w4787 , w2587 );
nor ( w4789 , w4788 , w2575 );
and ( w4790 , w4789 , w6110 );
not ( w4791 , w4790 );
and ( w4792 , w3154 , w4791 );
and ( w4793 , w2890 , w2883 );
and ( w4794 , w4793 , w4790 );
and ( w4795 , w4794 , w12142 );
not ( w4796 , w4795 );
and ( w4797 , w4796 , w3151 );
not ( w4798 , w4797 );
and ( w4799 , w4798 , w3615 );
not ( w4800 , w4799 );
and ( w4801 , w4800 , w310 );
and ( w4802 , w4801 , w11852 );
and ( w4803 , w4802 , w377 );
nor ( w4804 , w4803 , w2906 );
and ( w4805 , w4804 , w2908 );
nor ( w4806 , w4805 , w255 );
and ( w4807 , w377 , w4806 );
and ( w4808 , w19 , w11852 );
not ( w4809 , w4808 );
and ( w4810 , w4809 , g31 );
and ( w4811 , w4810 , w11852 );
and ( w4812 , w4811 , w310 );
not ( w4813 , w4812 );
and ( w4814 , w4813 , w3605 );
and ( w4815 , w4717 , w12144 );
and ( w4816 , w4815 , w12142 );
nor ( w4817 , w20 , w4816 );
and ( w4818 , w4817 , w5968 );
not ( w4819 , w4818 );
and ( w4820 , w4819 , w2582 );
not ( w4821 , w4820 );
and ( w4822 , w4821 , w2624 );
and ( w4823 , w4822 , w2587 );
nor ( w4824 , w4823 , w2575 );
and ( w4825 , w4824 , w6110 );
nor ( w4826 , w4814 , w4825 );
and ( w4827 , w4826 , g32 );
and ( w4828 , w4827 , g33 );
nor ( w4829 , w4825 , w4672 );
and ( w4830 , w11166 , w4829 );
and ( w4831 , w4830 , w4950 );
not ( w4832 , w4831 );
and ( w4833 , w4832 , w2582 );
not ( w4834 , w4833 );
and ( w4835 , w4834 , w2624 );
and ( w4836 , w4835 , w2587 );
nor ( w4837 , w4836 , w2575 );
and ( w4838 , w4837 , w6110 );
not ( w4839 , w4828 );
and ( w4840 , w4839 , w4838 );
nor ( w4841 , w4840 , w377 );
and ( w4842 , w11166 , w4841 );
and ( w4843 , w4842 , w4950 );
and ( w4844 , w4843 , w5898 );
and ( w4845 , w4844 , w11166 );
and ( w4846 , w4845 , w5968 );
not ( w4847 , w4846 );
and ( w4848 , w4847 , w2582 );
not ( w4849 , w4848 );
and ( w4850 , w4849 , w2624 );
and ( w4851 , w4850 , w2587 );
nor ( w4852 , w4851 , w2575 );
and ( w4853 , w4852 , w6110 );
and ( w4854 , w4853 , w2582 );
not ( w4855 , w4854 );
and ( w4856 , w4855 , w2587 );
nor ( w4857 , w4856 , w2575 );
and ( w4858 , w4857 , w6110 );
not ( w4859 , w4807 );
and ( w4860 , w4859 , w4858 );
nor ( w4861 , w20 , w4860 );
and ( w4862 , w4861 , w4950 );
and ( w4863 , w4862 , w5898 );
and ( w4864 , w4863 , w11166 );
and ( w4865 , w4864 , w12532 );
and ( w4866 , w4865 , w5968 );
not ( w4867 , w4866 );
and ( w4868 , w4867 , w2582 );
not ( w4869 , w4868 );
and ( w4870 , w4869 , w2624 );
and ( w4871 , w4870 , w2587 );
nor ( w4872 , w4871 , w2575 );
and ( w4873 , w4872 , w6110 );
not ( w4874 , w4792 );
and ( w4875 , w4874 , w4873 );
and ( w4876 , w4875 , w3615 );
not ( w4877 , w4876 );
and ( w4878 , w4877 , w310 );
and ( w4879 , w4878 , w11852 );
and ( w4880 , w4879 , w377 );
nor ( w4881 , w4880 , w2906 );
and ( w4882 , w4881 , w2908 );
nor ( w4883 , w4882 , w255 );
and ( w4884 , w377 , w4883 );
not ( w4885 , w4884 );
and ( w4886 , w4885 , w4858 );
nor ( w4887 , w4886 , w4617 );
and ( w4888 , w4887 , w5898 );
and ( w4889 , w4888 , w11166 );
and ( w4890 , w4889 , w12532 );
and ( w4891 , w4890 , w5968 );
not ( w4892 , w4891 );
and ( w4893 , w4892 , w2582 );
not ( w4894 , w4893 );
and ( w4895 , w4894 , w2587 );
nor ( w4896 , w4895 , w2575 );
and ( w4897 , w4896 , w6110 );
and ( w4898 , w4766 , w4897 );
nor ( w4899 , w20 , w4898 );
and ( w4900 , w4899 , w4950 );
and ( w4901 , w4900 , w5898 );
and ( w4902 , w4901 , w11166 );
and ( w4903 , w4902 , w12532 );
and ( w4904 , w4903 , w5968 );
not ( w4905 , w4904 );
and ( w4906 , w4905 , w2582 );
not ( w4907 , w4906 );
and ( w4908 , w4907 , w2624 );
and ( w4909 , w4908 , w2587 );
nor ( w4910 , w4909 , w2575 );
and ( w4911 , w4910 , w6110 );
not ( w4912 , w4760 );
and ( w4913 , w4912 , w4911 );
nor ( w4914 , w20 , w4913 );
and ( w4915 , w4914 , w4950 );
and ( w4916 , w4915 , w5898 );
and ( w4917 , w4916 , w11166 );
and ( w4918 , w4917 , w12532 );
and ( w4919 , w4918 , w5968 );
not ( w4920 , w4919 );
and ( w4921 , w4920 , w2582 );
not ( w4922 , w4921 );
and ( w4923 , w4922 , w2624 );
and ( w4924 , w4923 , w2587 );
nor ( w4925 , w4924 , w2575 );
and ( w4926 , w4925 , w6110 );
nor ( w4927 , w4660 , w4926 );
and ( w4928 , w4927 , w11852 );
and ( w4929 , w4928 , w8848 );
and ( w4930 , w4929 , w485 );
not ( w4931 , w4930 );
and ( w4932 , w4931 , w4911 );
nor ( w4933 , w4932 , w105 );
and ( w4934 , w4933 , w12532 );
and ( w4935 , w4934 , w5968 );
not ( w4936 , w4935 );
and ( w4937 , w4936 , w2582 );
not ( w4938 , w4937 );
and ( w4939 , w4938 , w2587 );
nor ( w4940 , w4939 , w2575 );
and ( w4941 , w4940 , w6110 );
not ( w4942 , w4690 );
and ( w4943 , w4942 , w4941 );
nor ( w4944 , w4943 , w19 );
and ( w4945 , w4944 , w485 );
not ( w4946 , w4945 );
and ( w4947 , w4946 , w4911 );
nor ( w4948 , w20 , w4947 );
and ( w4949 , w11166 , w4948 );
not ( w4950 , w4617 );
and ( w4951 , w4949 , w4950 );
and ( w4952 , w4951 , w5898 );
and ( w4953 , w4952 , w11166 );
and ( w4954 , w4953 , w5968 );
not ( w4955 , w4954 );
and ( w4956 , w4955 , w2582 );
not ( w4957 , w4956 );
and ( w4958 , w4957 , w2624 );
and ( w4959 , w4958 , w2587 );
nor ( w4960 , w4959 , w2575 );
and ( w4961 , w4960 , w6110 );
not ( w4962 , w4676 );
and ( w4963 , w4962 , w4961 );
nor ( w4964 , w4963 , w2994 );
and ( w4965 , w4964 , w11166 );
and ( w4966 , w4965 , w12532 );
and ( w4967 , w4966 , w5968 );
not ( w4968 , w4967 );
and ( w4969 , w4968 , w2582 );
not ( w4970 , w4969 );
and ( w4971 , w4970 , w2624 );
and ( w4972 , w4971 , w2587 );
nor ( w4973 , w4972 , w2575 );
and ( w4974 , w4973 , w6110 );
and ( w4975 , w4649 , w4974 );
not ( w4976 , w4975 );
and ( w4977 , w20 , w4976 );
not ( w4978 , w4977 );
and ( w4979 , w4978 , w4961 );
nor ( w4980 , w4979 , w2994 );
and ( w4981 , w4980 , w11166 );
and ( w4982 , w4981 , w12532 );
and ( w4983 , w4982 , w5968 );
not ( w4984 , w4983 );
and ( w4985 , w4984 , w2582 );
not ( w4986 , w4985 );
and ( w4987 , w4986 , w2624 );
and ( w4988 , w4987 , w2587 );
nor ( w4989 , w4988 , w2575 );
and ( w4990 , w4989 , w6110 );
not ( w4991 , w4990 );
and ( w4992 , w4991 , w312 );
not ( w4993 , w4992 );
and ( w4994 , w4993 , w4974 );
nor ( w4995 , w4994 , w2735 );
not ( w4996 , w4995 );
and ( w4997 , w4996 , w2582 );
not ( w4998 , w4997 );
and ( w4999 , w4998 , w2587 );
nor ( w5000 , w4999 , w2575 );
and ( w5001 , w3146 , w5000 );
nor ( w5002 , w5001 , w2735 );
not ( w5003 , w5002 );
and ( w5004 , w5003 , w2582 );
not ( w5005 , w5004 );
and ( w5006 , w5005 , w2624 );
and ( w5007 , w5006 , w2587 );
nor ( w5008 , w5007 , w2575 );
and ( w5009 , w5008 , w6110 );
not ( w5010 , w2980 );
and ( w5011 , w5010 , w5009 );
nor ( w5012 , w5011 , w384 );
and ( w5013 , w5012 , w12037 );
not ( w5014 , w5013 );
and ( w5015 , w5014 , w5000 );
nor ( w5016 , w5015 , w2735 );
not ( w5017 , w5016 );
and ( w5018 , w5017 , w2582 );
not ( w5019 , w5018 );
and ( w5020 , w5019 , w2624 );
and ( w5021 , w5020 , w2587 );
nor ( w5022 , w5021 , w2575 );
and ( w5023 , w5022 , w6110 );
nor ( w5024 , w2777 , w5023 );
and ( w5025 , w12921 , w5024 );
and ( w5026 , w5025 , w5968 );
not ( w5027 , w5026 );
and ( w5028 , w5027 , w2582 );
not ( w5029 , w5028 );
and ( w5030 , w5029 , w2624 );
and ( w5031 , w5030 , w2587 );
nor ( w5032 , w5031 , w2575 );
and ( w5033 , w5032 , w6110 );
not ( w5034 , w2717 );
and ( w5035 , w5034 , w5033 );
not ( w5036 , w5035 );
and ( w5037 , w5036 , w310 );
and ( w5038 , w5037 , w11852 );
and ( w5039 , w5038 , w12532 );
nor ( w5040 , w5039 , w2906 );
and ( w5041 , w5040 , w2908 );
not ( w5042 , w5041 );
and ( w5043 , w5042 , w377 );
not ( w5044 , w5043 );
and ( w5045 , w5044 , w2971 );
and ( w5046 , w5045 , w8363 );
nor ( w5047 , w5046 , w2883 );
not ( w5048 , w2888 );
and ( w5049 , w5047 , w5048 );
and ( w5050 , w5049 , w8363 );
and ( w5051 , w5050 , w12144 );
and ( w5052 , w5051 , w239 );
not ( w5053 , w5052 );
and ( w5054 , w5053 , w3005 );
and ( w5055 , w5054 , w2976 );
and ( w5056 , w5055 , w11166 );
nor ( w5057 , w5056 , w18 );
and ( w5058 , w5057 , w11166 );
not ( w5059 , w4677 );
and ( w5060 , w5059 , w3097 );
not ( w5061 , w5033 );
and ( w5062 , w5061 , w310 );
and ( w5063 , w5062 , w11852 );
and ( w5064 , w5063 , w12532 );
and ( w5065 , w5064 , w377 );
not ( w5066 , w5065 );
and ( w5067 , w5066 , w2775 );
and ( w5068 , w5067 , w2664 );
not ( w5069 , w3899 );
and ( w5070 , w5069 , w2713 );
not ( w5071 , w5070 );
and ( w5072 , w5071 , w255 );
nor ( w5073 , w5072 , w43 );
and ( w5074 , w5073 , w4393 );
nor ( w5075 , w5074 , w43 );
and ( w5076 , w5075 , w5370 );
nor ( w5077 , w5076 , w2592 );
and ( w5078 , w5077 , w2976 );
and ( w5079 , w5078 , w3124 );
nor ( w5080 , w5079 , w3116 );
nor ( w5081 , w5080 , w105 );
and ( w5082 , w5081 , w12498 );
and ( w5083 , w5082 , w2775 );
nor ( w5084 , w5083 , w2961 );
and ( w5085 , w5084 , w12498 );
not ( w5086 , w5085 );
and ( w5087 , w5086 , w3875 );
not ( w5088 , w5087 );
and ( w5089 , w5088 , g33 );
and ( w5090 , w5089 , g32 );
not ( w5091 , w5090 );
and ( w5092 , w5091 , g32 );
and ( w5093 , w5092 , g33 );
not ( w5094 , w2649 );
and ( w5095 , w5093 , w5094 );
not ( w5096 , w5095 );
and ( w5097 , w5096 , w312 );
and ( w5098 , w5097 , w12717 );
and ( w5099 , w5098 , w384 );
and ( w5100 , w12921 , w5099 );
not ( w5101 , w2582 );
and ( w5102 , w5101 , w2624 );
and ( w5103 , w5102 , w2587 );
nor ( w5104 , w5103 , w2575 );
and ( w5105 , w5104 , w6110 );
not ( w5106 , w5100 );
and ( w5107 , w5106 , w5105 );
nor ( w5108 , w5107 , w2735 );
not ( w5109 , w5108 );
and ( w5110 , w5109 , w2582 );
not ( w5111 , w5110 );
and ( w5112 , w5111 , w2624 );
and ( w5113 , w5112 , w2587 );
nor ( w5114 , w5113 , w2575 );
and ( w5115 , w5114 , w6110 );
and ( w5116 , w5068 , w5115 );
and ( w5117 , w5116 , w5105 );
and ( w5118 , w5117 , w5000 );
nor ( w5119 , w5118 , w2735 );
not ( w5120 , w5119 );
and ( w5121 , w5120 , w2582 );
not ( w5122 , w5121 );
and ( w5123 , w5122 , w2587 );
nor ( w5124 , w5123 , w2575 );
and ( w5125 , w5124 , w6110 );
and ( w5126 , w5060 , w5125 );
nor ( w5127 , w5126 , g29 );
not ( w5128 , w5127 );
and ( w5129 , w5128 , w2775 );
and ( w5130 , w5129 , w2664 );
and ( w5131 , w5130 , w5105 );
and ( w5132 , w5131 , w5000 );
and ( w5133 , w5132 , w2582 );
not ( w5134 , w5133 );
and ( w5135 , w5134 , w2587 );
nor ( w5136 , w5135 , w2575 );
and ( w5137 , w5136 , w6110 );
not ( w5138 , w5058 );
and ( w5139 , w5138 , w5137 );
and ( w5140 , w5139 , w5115 );
nor ( w5141 , w20 , w5140 );
not ( w5142 , w5141 );
and ( w5143 , w5142 , w5105 );
and ( w5144 , w5143 , w5000 );
nor ( w5145 , w5144 , w2735 );
not ( w5146 , w5145 );
and ( w5147 , w5146 , w2582 );
not ( w5148 , w5147 );
and ( w5149 , w5148 , w2624 );
and ( w5150 , w5149 , w2587 );
nor ( w5151 , w5150 , w2575 );
and ( w5152 , w5151 , w6110 );
not ( w5153 , w2653 );
and ( w5154 , w5153 , w5152 );
nor ( w5155 , w5154 , g29 );
and ( w5156 , w5155 , w3867 );
and ( w5157 , w5156 , w377 );
not ( w5158 , w5157 );
and ( w5159 , w5158 , w2971 );
nor ( w5160 , w35 , w5159 );
not ( w5161 , w5160 );
and ( w5162 , w5161 , w3005 );
and ( w5163 , w5162 , w2976 );
and ( w5164 , w5163 , w11166 );
not ( w5165 , w5164 );
and ( w5166 , w5165 , w4205 );
and ( w5167 , w5166 , w12919 );
and ( w5168 , w5167 , w11166 );
not ( w5169 , w5168 );
and ( w5170 , w5169 , w5137 );
and ( w5171 , w5170 , w5115 );
nor ( w5172 , w20 , w5171 );
not ( w5173 , w5172 );
and ( w5174 , w5173 , w5105 );
and ( w5175 , w5174 , w5000 );
nor ( w5176 , w5175 , w2735 );
not ( w5177 , w5176 );
and ( w5178 , w5177 , w2582 );
not ( w5179 , w5178 );
and ( w5180 , w5179 , w2624 );
and ( w5181 , w5180 , w2587 );
nor ( w5182 , w5181 , w2575 );
and ( w5183 , w5182 , w6110 );
and ( w5184 , w2593 , w5183 );
and ( w5185 , w5184 , w2582 );
not ( w5186 , w5185 );
and ( w5187 , w5186 , w2587 );
nor ( w5188 , w5187 , w2575 );
and ( w5189 , w5188 , w6110 );
and ( w5190 , w5189 , w19 );
and ( w5191 , w5190 , w5183 );
and ( w5192 , w5191 , w2582 );
not ( w5193 , w5192 );
and ( w5194 , w5193 , w2624 );
and ( w5195 , w5194 , w2587 );
nor ( w5196 , w5195 , w2575 );
and ( w5197 , w5196 , w19 );
and ( w5198 , w5197 , w12080 );
nor ( w5199 , w5198 , w2994 );
and ( w5200 , w20 , w5199 );
not ( w5201 , w5200 );
and ( w5202 , w5201 , w5105 );
nor ( w5203 , w384 , w308 );
nor ( w5204 , w5203 , w310 );
and ( w5205 , w5204 , w384 );
nor ( w5206 , w5205 , w308 );
nor ( w5207 , w3734 , w2888 );
nor ( w5208 , w5207 , w48 );
nor ( w5209 , w5208 , w2961 );
and ( w5210 , w5209 , w12498 );
and ( w5211 , w377 , w12080 );
and ( w5212 , w5211 , w2587 );
nor ( w5213 , w5210 , w5212 );
and ( w5214 , w5874 , w20 );
and ( w5215 , w5214 , w11166 );
and ( w5216 , w20 , w5215 );
and ( w5217 , w5216 , w12717 );
nor ( w5218 , w2888 , w3744 );
and ( w5219 , w5218 , w8848 );
and ( w5220 , w5219 , w5898 );
nor ( w5221 , w5220 , w377 );
and ( w5222 , w2971 , w3017 );
and ( w5223 , w5222 , w2976 );
nor ( w5224 , w5223 , w18 );
not ( w5225 , w5224 );
and ( w5226 , w5225 , w2775 );
nor ( w5227 , w20 , w5226 );
and ( w5228 , w5227 , w5968 );
not ( w5229 , w5228 );
and ( w5230 , w5229 , w2582 );
not ( w5231 , w5230 );
and ( w5232 , w5231 , w2624 );
and ( w5233 , w5232 , w2587 );
nor ( w5234 , w5233 , w2575 );
and ( w5235 , w5234 , w6110 );
and ( w5236 , w5221 , w5235 );
and ( w5237 , w5236 , w2775 );
nor ( w5238 , w5237 , w2961 );
nor ( w5239 , w377 , w5238 );
nor ( w5240 , w20 , w5239 );
and ( w5241 , w5240 , w5968 );
not ( w5242 , w5241 );
and ( w5243 , w5242 , w2582 );
not ( w5244 , w5243 );
and ( w5245 , w5244 , w2624 );
and ( w5246 , w5245 , w2587 );
nor ( w5247 , w5246 , w2575 );
and ( w5248 , w5247 , w6110 );
and ( w5249 , w11852 , w5248 );
nor ( w5250 , w5249 , w5203 );
nor ( w5251 , w5250 , w19 );
nor ( w5252 , w19 , w105 );
and ( w5253 , w5252 , w5968 );
and ( w5254 , w5253 , w2624 );
and ( w5255 , w5254 , w2587 );
nor ( w5256 , w5255 , w2575 );
and ( w5257 , w377 , w5727 );
nor ( w5258 , w377 , w5235 );
not ( w5259 , w5258 );
and ( w5260 , w5259 , w5183 );
and ( w5261 , w5260 , w2582 );
not ( w5262 , w5261 );
and ( w5263 , w5262 , w2587 );
nor ( w5264 , w5263 , w2575 );
and ( w5265 , w5264 , w6110 );
and ( w5266 , w19 , w2593 );
nor ( w5267 , w5218 , w377 );
nor ( w5268 , w5267 , w3696 );
not ( w5269 , w5268 );
and ( w5270 , w5269 , w2775 );
and ( w5271 , w12498 , w5270 );
nor ( w5272 , w5271 , w310 );
and ( w5273 , w12921 , w5272 );
and ( w5274 , w5273 , w12037 );
not ( w5275 , w5274 );
and ( w5276 , w5275 , w5183 );
nor ( w5277 , w5276 , w2735 );
not ( w5278 , w5277 );
and ( w5279 , w5278 , w2582 );
not ( w5280 , w5279 );
and ( w5281 , w5280 , w2624 );
and ( w5282 , w5281 , w2587 );
nor ( w5283 , w5282 , w2575 );
and ( w5284 , w5283 , w6110 );
nor ( w5285 , w5266 , w5284 );
and ( w5286 , w377 , w5285 );
nor ( w5287 , w4786 , w3744 );
and ( w5288 , w5287 , w5364 );
and ( w5289 , w5288 , w8848 );
not ( w5290 , w5289 );
and ( w5291 , w5290 , w2976 );
nor ( w5292 , w5291 , w2961 );
and ( w5293 , w5292 , w5597 );
not ( w5294 , w5293 );
and ( w5295 , w5294 , w3106 );
nor ( w5296 , w5295 , w310 );
and ( w5297 , w5296 , w12037 );
not ( w5298 , w5297 );
and ( w5299 , w5298 , w5183 );
nor ( w5300 , w5299 , w2735 );
not ( w5301 , w5300 );
and ( w5302 , w5301 , w2582 );
not ( w5303 , w5302 );
and ( w5304 , w5303 , w2587 );
nor ( w5305 , w5304 , w2575 );
and ( w5306 , w5305 , w6110 );
nor ( w5307 , w19 , w5306 );
and ( w5308 , w5307 , w12717 );
and ( w5309 , w5308 , w12037 );
not ( w5310 , w5309 );
and ( w5311 , w5310 , w5183 );
nor ( w5312 , w5311 , w2735 );
not ( w5313 , w5312 );
and ( w5314 , w5313 , w2582 );
not ( w5315 , w5314 );
and ( w5316 , w5315 , w2587 );
nor ( w5317 , w5316 , w2575 );
not ( w5318 , w5286 );
and ( w5319 , w5318 , w5317 );
and ( w5320 , w5319 , w11166 );
and ( w5321 , w4243 , w2961 );
and ( w5322 , w5321 , w5183 );
nor ( w5323 , w5322 , w2735 );
not ( w5324 , w5323 );
and ( w5325 , w5324 , w2582 );
not ( w5326 , w5325 );
and ( w5327 , w5326 , w2587 );
nor ( w5328 , w5327 , w2575 );
nor ( w5329 , w5320 , w5328 );
and ( w5330 , w5329 , w5898 );
and ( w5331 , w5330 , w48 );
nor ( w5332 , w5331 , w2592 );
not ( w5333 , w3683 );
and ( w5334 , w5218 , w5333 );
and ( w5335 , w5334 , w5366 );
and ( w5336 , w5335 , w11140 );
and ( w5337 , w5336 , w5422 );
and ( w5338 , w5337 , w5370 );
and ( w5339 , w5338 , w8848 );
not ( w5340 , w5339 );
and ( w5341 , w5340 , w2976 );
nor ( w5342 , w5341 , w2961 );
and ( w5343 , w5342 , w5597 );
not ( w5344 , w5343 );
and ( w5345 , w5344 , w3106 );
and ( w5346 , w5345 , w12144 );
nor ( w5347 , w20 , w5346 );
and ( w5348 , w5347 , w5968 );
not ( w5349 , w5348 );
and ( w5350 , w5349 , w2582 );
not ( w5351 , w5350 );
and ( w5352 , w5351 , w2624 );
and ( w5353 , w5352 , w2587 );
nor ( w5354 , w5353 , w2575 );
and ( w5355 , w5354 , w6110 );
and ( w5356 , w12498 , w5355 );
and ( w5357 , w5207 , w8848 );
and ( w5358 , w5357 , w12919 );
not ( w5359 , w5358 );
and ( w5360 , w5359 , w2593 );
and ( w5361 , w5360 , w4218 );
nor ( w5362 , w5361 , w5328 );
and ( w5363 , w377 , w5362 );
not ( w5364 , w3689 );
and ( w5365 , w5218 , w5364 );
not ( w5366 , w3233 );
and ( w5367 , w5365 , w5366 );
and ( w5368 , w5367 , w11140 );
and ( w5369 , w5368 , w5422 );
not ( w5370 , w2680 );
and ( w5371 , w5369 , w5370 );
not ( w5372 , w5371 );
and ( w5373 , w5372 , w2976 );
nor ( w5374 , w5373 , w2961 );
and ( w5375 , w5374 , w12498 );
and ( w5376 , w5375 , w5597 );
not ( w5377 , w5376 );
and ( w5378 , w5377 , w3106 );
and ( w5379 , w5378 , w12144 );
nor ( w5380 , w20 , w5379 );
and ( w5381 , w5380 , w5968 );
and ( w5382 , w5381 , w2624 );
and ( w5383 , w5382 , w2587 );
nor ( w5384 , w5383 , w2575 );
and ( w5385 , w5384 , w6110 );
not ( w5386 , w5363 );
and ( w5387 , w5386 , w5385 );
nor ( w5388 , w5387 , w5284 );
and ( w5389 , w5388 , w12080 );
and ( w5390 , w5389 , w12717 );
and ( w5391 , w11852 , w5390 );
and ( w5392 , w12921 , w5391 );
and ( w5393 , w5392 , w12037 );
not ( w5394 , w5393 );
and ( w5395 , w5394 , w5183 );
nor ( w5396 , w5395 , w2735 );
not ( w5397 , w5396 );
and ( w5398 , w5397 , w2582 );
not ( w5399 , w5398 );
and ( w5400 , w5399 , w2624 );
and ( w5401 , w5400 , w2587 );
nor ( w5402 , w5401 , w2575 );
and ( w5403 , w5402 , w6110 );
nor ( w5404 , w5356 , w5403 );
and ( w5405 , w5404 , w12144 );
and ( w5406 , w12498 , w5306 );
nor ( w5407 , w5406 , w5284 );
and ( w5408 , w39 , w12144 );
nor ( w5409 , w5408 , w45 );
and ( w5410 , w5409 , w11347 );
and ( w5411 , w5410 , w37 );
and ( w5412 , w5411 , w8848 );
not ( w5413 , w5412 );
and ( w5414 , w5413 , w2976 );
nor ( w5415 , w5414 , w2961 );
and ( w5416 , w5415 , w12498 );
nor ( w5417 , w2883 , w2888 );
and ( w5418 , w5417 , w239 );
and ( w5419 , w5418 , w11347 );
and ( w5420 , w7803 , w5419 );
and ( w5421 , w5420 , w11140 );
not ( w5422 , w2674 );
and ( w5423 , w5421 , w5422 );
and ( w5424 , w235 , w5968 );
and ( w5425 , w5424 , w2587 );
nor ( w5426 , w5425 , w2575 );
and ( w5427 , w5426 , w6110 );
not ( w5428 , w5423 );
and ( w5429 , w5428 , w5427 );
and ( w5430 , w5429 , w12144 );
nor ( w5431 , w5430 , w45 );
and ( w5432 , w5431 , w8848 );
not ( w5433 , w5432 );
and ( w5434 , w5433 , w2976 );
nor ( w5435 , w5434 , w2961 );
and ( w5436 , w5435 , w12498 );
and ( w5437 , w5436 , w5597 );
not ( w5438 , w5437 );
and ( w5439 , w5438 , w3106 );
nor ( w5440 , w37 , w5439 );
and ( w5441 , w5440 , w12717 );
and ( w5442 , w12921 , w5441 );
and ( w5443 , w5442 , w5968 );
not ( w5444 , w5443 );
and ( w5445 , w5444 , w2582 );
not ( w5446 , w5445 );
and ( w5447 , w5446 , w2624 );
and ( w5448 , w5447 , w2587 );
nor ( w5449 , w5448 , w2575 );
and ( w5450 , w5449 , w6110 );
not ( w5451 , w5416 );
and ( w5452 , w5451 , w5450 );
nor ( w5453 , w5452 , w3116 );
not ( w5454 , w5453 );
and ( w5455 , w5454 , w3106 );
nor ( w5456 , w3734 , w4786 );
and ( w5457 , w5456 , w8848 );
not ( w5458 , w5457 );
and ( w5459 , w5458 , w2593 );
nor ( w5460 , w5459 , w18 );
not ( w5461 , w5460 );
and ( w5462 , w5461 , w4218 );
nor ( w5463 , w5462 , w5328 );
and ( w5464 , w377 , w5463 );
and ( w5465 , w5464 , w12080 );
and ( w5466 , w5465 , w12717 );
and ( w5467 , w11852 , w5466 );
and ( w5468 , w12921 , w5467 );
not ( w5469 , w5468 );
and ( w5470 , w5469 , w5183 );
nor ( w5471 , w5470 , w2735 );
not ( w5472 , w5471 );
and ( w5473 , w5472 , w2582 );
not ( w5474 , w5473 );
and ( w5475 , w5474 , w2624 );
and ( w5476 , w5475 , w2587 );
nor ( w5477 , w5476 , w2575 );
and ( w5478 , w5477 , w6110 );
and ( w5479 , w5455 , w5478 );
nor ( w5480 , w5479 , w255 );
and ( w5481 , w5480 , w12717 );
and ( w5482 , w12921 , w5481 );
and ( w5483 , w5482 , w5968 );
not ( w5484 , w5483 );
and ( w5485 , w5484 , w2582 );
not ( w5486 , w5485 );
and ( w5487 , w5486 , w2624 );
and ( w5488 , w5487 , w2587 );
nor ( w5489 , w5488 , w2575 );
and ( w5490 , w5489 , w6110 );
not ( w5491 , w5490 );
and ( w5492 , w5407 , w5491 );
and ( w5493 , w5492 , w12080 );
and ( w5494 , w5493 , w12717 );
and ( w5495 , w5494 , w12037 );
not ( w5496 , w5495 );
and ( w5497 , w5496 , w5183 );
nor ( w5498 , w5497 , w2735 );
not ( w5499 , w5498 );
and ( w5500 , w5499 , w2582 );
not ( w5501 , w5500 );
and ( w5502 , w5501 , w2587 );
nor ( w5503 , w5502 , w2575 );
and ( w5504 , w5503 , w6110 );
not ( w5505 , w5405 );
and ( w5506 , w5505 , w5504 );
nor ( w5507 , w5506 , w48 );
and ( w5508 , w5507 , w12080 );
and ( w5509 , w5508 , w5968 );
not ( w5510 , w5509 );
and ( w5511 , w5510 , w2582 );
not ( w5512 , w5511 );
and ( w5513 , w5512 , w2587 );
nor ( w5514 , w5513 , w2575 );
and ( w5515 , w5514 , w6110 );
and ( w5516 , w5332 , w5515 );
nor ( w5517 , w5516 , w5248 );
and ( w5518 , w5517 , w12532 );
and ( w5519 , w5518 , w12080 );
and ( w5520 , w5519 , w12717 );
and ( w5521 , w11852 , w5520 );
and ( w5522 , w5521 , w12037 );
not ( w5523 , w5522 );
and ( w5524 , w5523 , w5183 );
nor ( w5525 , w5524 , w2735 );
not ( w5526 , w5525 );
and ( w5527 , w5526 , w2582 );
not ( w5528 , w5527 );
and ( w5529 , w5528 , w2624 );
and ( w5530 , w5529 , w2587 );
nor ( w5531 , w5530 , w2575 );
and ( w5532 , w5531 , w6110 );
and ( w5533 , w5265 , w5532 );
and ( w5534 , w5533 , w5183 );
and ( w5535 , w5534 , w2589 );
not ( w5536 , w789 );
and ( w5537 , w5535 , w5536 );
nor ( w5538 , w5537 , w377 );
not ( w5539 , w5538 );
and ( w5540 , w5539 , w19 );
and ( w5541 , w5540 , w5532 );
and ( w5542 , w5541 , w6110 );
and ( w5543 , w5542 , w5183 );
nor ( w5544 , w5543 , w2735 );
not ( w5545 , w5544 );
and ( w5546 , w5545 , w2582 );
not ( w5547 , w5546 );
and ( w5548 , w5547 , w2624 );
and ( w5549 , w5548 , w2587 );
nor ( w5550 , w5549 , w2575 );
and ( w5551 , w5550 , w6110 );
not ( w5552 , w5257 );
and ( w5553 , w5552 , w5551 );
nor ( w5554 , w5553 , w105 );
not ( w5555 , w5554 );
and ( w5556 , w5555 , w2976 );
nor ( w5557 , w5556 , w3113 );
not ( w5558 , w5557 );
and ( w5559 , w5558 , w3097 );
and ( w5560 , w5559 , w8640 );
nor ( w5561 , w20 , w5560 );
nor ( w5562 , w5561 , w2592 );
and ( w5563 , w5562 , w5183 );
nor ( w5564 , w5563 , w2735 );
not ( w5565 , w5564 );
and ( w5566 , w5565 , w2582 );
not ( w5567 , w5566 );
and ( w5568 , w5567 , w2624 );
and ( w5569 , w5568 , w2587 );
nor ( w5570 , w5569 , w2575 );
and ( w5571 , w5570 , w6110 );
nor ( w5572 , w5251 , w5571 );
not ( w5573 , w5572 );
and ( w5574 , w5573 , w5532 );
nor ( w5575 , w5574 , w310 );
and ( w5576 , w3433 , w3431 );
and ( w5577 , w5576 , w4200 );
and ( w5578 , w5577 , w2587 );
not ( w5579 , w5578 );
and ( w5580 , g31 , w5579 );
nor ( w5581 , w5580 , w310 );
and ( w5582 , w5581 , w2587 );
and ( w5583 , w3623 , w5582 );
and ( w5584 , w5583 , w12717 );
and ( w5585 , w5584 , w2587 );
not ( w5586 , w5585 );
and ( w5587 , w5586 , w255 );
nor ( w5588 , w5587 , w310 );
and ( w5589 , w5588 , w2587 );
and ( w5590 , w384 , w5589 );
nor ( w5591 , w5590 , w789 );
and ( w5592 , w2674 , w12144 );
and ( w5593 , w5592 , w12142 );
and ( w5594 , w5593 , w12921 );
and ( w5595 , w5594 , w2976 );
nor ( w5596 , w5595 , w20 );
not ( w5597 , w3116 );
and ( w5598 , w5596 , w5597 );
not ( w5599 , w5598 );
and ( w5600 , w5599 , w2775 );
and ( w5601 , w12498 , w5600 );
nor ( w5602 , w5601 , w2735 );
not ( w5603 , w5602 );
and ( w5604 , w5603 , w2582 );
not ( w5605 , w5604 );
and ( w5606 , w5605 , w2624 );
and ( w5607 , w5606 , w2587 );
nor ( w5608 , w5607 , w2575 );
and ( w5609 , w5608 , w6110 );
and ( w5610 , w12921 , w5609 );
nor ( w5611 , w5610 , w2735 );
and ( w5612 , w5611 , w2624 );
and ( w5613 , w5612 , w2587 );
nor ( w5614 , w5613 , w2575 );
and ( w5615 , w5614 , w6110 );
nor ( w5616 , w5615 , w5196 );
and ( w5617 , w5616 , w5898 );
and ( w5618 , w5617 , w20 );
and ( w5619 , w5618 , w11166 );
and ( w5620 , w20 , w5619 );
not ( w5621 , w5620 );
and ( w5622 , w5621 , w5105 );
and ( w5623 , w3734 , w12142 );
nor ( w5624 , w5623 , w2888 );
and ( w5625 , w5624 , w12919 );
and ( w5626 , w5625 , w11166 );
and ( w5627 , w12921 , w5626 );
and ( w5628 , w2664 , w2582 );
not ( w5629 , w5628 );
and ( w5630 , w5629 , w2587 );
nor ( w5631 , w5630 , w2575 );
and ( w5632 , w5631 , w6110 );
and ( w5633 , w2664 , w5632 );
and ( w5634 , w5633 , w2582 );
not ( w5635 , w5634 );
and ( w5636 , w5635 , w2587 );
nor ( w5637 , w5636 , w2575 );
and ( w5638 , w5637 , w6110 );
not ( w5639 , w5627 );
and ( w5640 , w5639 , w5638 );
nor ( w5641 , w5640 , w2735 );
not ( w5642 , w5641 );
and ( w5643 , w5642 , w2582 );
not ( w5644 , w5643 );
and ( w5645 , w5644 , w2624 );
and ( w5646 , w5645 , w2587 );
nor ( w5647 , w5646 , w2575 );
and ( w5648 , w5647 , w6110 );
not ( w5649 , w4200 );
and ( w5650 , w5648 , w5649 );
not ( w5651 , w5650 );
and ( w5652 , w384 , w5651 );
not ( w5653 , w5571 );
and ( w5654 , w5652 , w5653 );
not ( w5655 , w5654 );
and ( w5656 , w5655 , w5532 );
nor ( w5657 , w5656 , w310 );
nor ( w5658 , w5657 , w308 );
and ( w5659 , w5898 , w20 );
and ( w5660 , w5659 , w11166 );
and ( w5661 , w20 , w5660 );
not ( w5662 , w5661 );
and ( w5663 , w5662 , w5105 );
and ( w5664 , w5663 , w5648 );
and ( w5665 , w19 , w5105 );
not ( w5666 , w5665 );
and ( w5667 , w5666 , w20 );
and ( w5668 , w2713 , w3005 );
not ( w5669 , w2906 );
and ( w5670 , w5668 , w5669 );
and ( w5671 , w5670 , w2908 );
not ( w5672 , w5671 );
and ( w5673 , w5672 , w377 );
and ( w5674 , w5235 , w5183 );
and ( w5675 , w5674 , w2582 );
not ( w5676 , w5675 );
and ( w5677 , w5676 , w2587 );
nor ( w5678 , w5677 , w2575 );
not ( w5679 , w5673 );
and ( w5680 , w5679 , w5678 );
and ( w5681 , w5680 , w8640 );
and ( w5682 , w5681 , w19 );
and ( w5683 , w5682 , w2976 );
and ( w5684 , w5683 , w11166 );
nor ( w5685 , w5684 , w18 );
and ( w5686 , w5685 , w11166 );
not ( w5687 , w5686 );
and ( w5688 , w5687 , w5638 );
nor ( w5689 , w20 , w5688 );
not ( w5690 , w5689 );
and ( w5691 , w5690 , w5183 );
nor ( w5692 , w5691 , w2735 );
not ( w5693 , w5692 );
and ( w5694 , w5693 , w2582 );
not ( w5695 , w5694 );
and ( w5696 , w5695 , w2624 );
and ( w5697 , w5696 , w2587 );
nor ( w5698 , w5697 , w2575 );
and ( w5699 , w5698 , w6110 );
not ( w5700 , w5667 );
and ( w5701 , w5700 , w5699 );
and ( w5702 , w5701 , w5183 );
nor ( w5703 , w5702 , w2735 );
not ( w5704 , w5703 );
and ( w5705 , w5704 , w2582 );
not ( w5706 , w5705 );
and ( w5707 , w5706 , w2587 );
nor ( w5708 , w5707 , w2575 );
and ( w5709 , w5708 , w6110 );
nor ( w5710 , w5664 , w5709 );
and ( w5711 , w5710 , w310 );
nor ( w5712 , w5711 , w2592 );
nor ( w5713 , w5712 , w384 );
and ( w5714 , w310 , w5713 );
and ( w5715 , w4677 , w12080 );
not ( w5716 , w5715 );
and ( w5717 , w5716 , w3116 );
and ( w5718 , w5717 , w3113 );
and ( w5719 , w5718 , w18 );
and ( w5720 , w5719 , w12921 );
and ( w5721 , w5720 , w2994 );
nor ( w5722 , w3734 , w2883 );
nor ( w5723 , w5722 , w20 );
and ( w5724 , w5723 , w12142 );
and ( w5725 , w12921 , w5724 );
nor ( w5726 , w5725 , w105 );
not ( w5727 , w5256 );
and ( w5728 , w5726 , w5727 );
and ( w5729 , w3098 , w2582 );
not ( w5730 , w5729 );
and ( w5731 , w5730 , w2587 );
nor ( w5732 , w5731 , w2575 );
and ( w5733 , w5732 , w6110 );
and ( w5734 , w5733 , w2582 );
not ( w5735 , w5734 );
and ( w5736 , w5735 , w2624 );
and ( w5737 , w5736 , w2587 );
nor ( w5738 , w5737 , w2575 );
and ( w5739 , w5738 , w6110 );
not ( w5740 , w5728 );
and ( w5741 , w5740 , w5739 );
and ( w5742 , w5741 , w377 );
and ( w5743 , w12921 , w2883 );
and ( w5744 , w5743 , w3106 );
and ( w5745 , w12921 , w5744 );
and ( w5746 , w5745 , w2888 );
nor ( w5747 , w5746 , w3744 );
not ( w5748 , w3696 );
and ( w5749 , w5747 , w5748 );
not ( w5750 , w5615 );
and ( w5751 , w5749 , w5750 );
nor ( w5752 , w5751 , w377 );
nor ( w5753 , w5752 , w2961 );
nor ( w5754 , w377 , w5753 );
nor ( w5755 , w5754 , w2735 );
and ( w5756 , w5755 , w2624 );
and ( w5757 , w5756 , w2587 );
nor ( w5758 , w5757 , w2575 );
nor ( w5759 , w5742 , w5758 );
nor ( w5760 , w5759 , w3431 );
and ( w5761 , w12080 , w5760 );
and ( w5762 , w5749 , w5589 );
nor ( w5763 , w2575 , w2592 );
and ( w5764 , w5763 , w5265 );
and ( w5765 , w5764 , w8640 );
and ( w5766 , w5765 , w19 );
and ( w5767 , w5766 , w11166 );
and ( w5768 , w5767 , w12498 );
nor ( w5769 , w5768 , w2961 );
and ( w5770 , w5769 , w12498 );
nor ( w5771 , w5770 , w2592 );
and ( w5772 , w5771 , w5183 );
nor ( w5773 , w5772 , w2735 );
not ( w5774 , w5773 );
and ( w5775 , w5774 , w2582 );
not ( w5776 , w5775 );
and ( w5777 , w5776 , w2624 );
and ( w5778 , w5777 , w2587 );
nor ( w5779 , w5778 , w2575 );
and ( w5780 , w5779 , w6110 );
not ( w5781 , w5780 );
and ( w5782 , w5762 , w5781 );
nor ( w5783 , w5782 , w789 );
and ( w5784 , w5783 , w2908 );
and ( w5785 , w5784 , w12498 );
nor ( w5786 , w5785 , w2961 );
nor ( w5787 , w377 , w5786 );
and ( w5788 , w5787 , w11226 );
and ( w5789 , w5788 , w13211 );
and ( w5790 , w5789 , w308 );
nor ( w5791 , w5790 , w312 );
not ( w5792 , w5791 );
and ( w5793 , w5792 , w5183 );
nor ( w5794 , w5793 , w2735 );
not ( w5795 , w5794 );
and ( w5796 , w5795 , w2582 );
not ( w5797 , w5796 );
and ( w5798 , w5797 , w2624 );
and ( w5799 , w5798 , w2587 );
nor ( w5800 , w5799 , w2575 );
and ( w5801 , w5800 , w6110 );
nor ( w5802 , w5761 , w5801 );
and ( w5803 , w5802 , w12717 );
not ( w5804 , w5803 );
and ( w5805 , w5804 , w308 );
and ( w5806 , w5805 , w6110 );
nor ( w5807 , w5806 , w312 );
not ( w5808 , w5807 );
and ( w5809 , w5808 , w5183 );
nor ( w5810 , w5809 , w2735 );
not ( w5811 , w5810 );
and ( w5812 , w5811 , w2582 );
not ( w5813 , w5812 );
and ( w5814 , w5813 , w2624 );
and ( w5815 , w5814 , w2587 );
nor ( w5816 , w5815 , w2575 );
and ( w5817 , w5816 , w6110 );
nor ( w5818 , w5721 , w5817 );
not ( w5819 , w5818 );
and ( w5820 , w5819 , w308 );
nor ( w5821 , w5820 , w312 );
not ( w5822 , w5821 );
and ( w5823 , w5822 , w5183 );
nor ( w5824 , w5823 , w2735 );
not ( w5825 , w5824 );
and ( w5826 , w5825 , w2582 );
not ( w5827 , w5826 );
and ( w5828 , w5827 , w2587 );
nor ( w5829 , w5828 , w2575 );
not ( w5830 , w5714 );
and ( w5831 , w5830 , w5829 );
and ( w5832 , w5831 , w11226 );
and ( w5833 , w5832 , w13211 );
and ( w5834 , w5833 , w308 );
nor ( w5835 , w5834 , w312 );
not ( w5836 , w5835 );
and ( w5837 , w5836 , w5183 );
nor ( w5838 , w5837 , w2735 );
not ( w5839 , w5838 );
and ( w5840 , w5839 , w2582 );
not ( w5841 , w5840 );
and ( w5842 , w5841 , w2624 );
and ( w5843 , w5842 , w2587 );
nor ( w5844 , w5843 , w2575 );
and ( w5845 , w5844 , w6110 );
nor ( w5846 , w5658 , w5845 );
and ( w5847 , w5846 , w12037 );
not ( w5848 , w5847 );
and ( w5849 , w5848 , w5183 );
nor ( w5850 , w5849 , w2735 );
not ( w5851 , w5850 );
and ( w5852 , w5851 , w2582 );
not ( w5853 , w5852 );
and ( w5854 , w5853 , w2587 );
nor ( w5855 , w5854 , w2575 );
and ( w5856 , w5855 , w6110 );
and ( w5857 , w5622 , w5856 );
nor ( w5858 , w5857 , w310 );
nor ( w5859 , w5858 , w308 );
nor ( w5860 , w5859 , w5845 );
and ( w5861 , w5860 , w12037 );
not ( w5862 , w5861 );
and ( w5863 , w5862 , w5183 );
nor ( w5864 , w5863 , w2735 );
not ( w5865 , w5864 );
and ( w5866 , w5865 , w2582 );
not ( w5867 , w5866 );
and ( w5868 , w5867 , w2624 );
and ( w5869 , w5868 , w2587 );
nor ( w5870 , w5869 , w2575 );
and ( w5871 , w5870 , w6110 );
nor ( w5872 , w5591 , w5871 );
and ( w5873 , w5872 , w12498 );
not ( w5874 , w5196 );
and ( w5875 , w5873 , w5874 );
and ( w5876 , w5875 , w5898 );
and ( w5877 , w5876 , w20 );
and ( w5878 , w5877 , w11166 );
and ( w5879 , w20 , w5878 );
not ( w5880 , w5879 );
and ( w5881 , w5880 , w5105 );
and ( w5882 , w5881 , w5856 );
and ( w5883 , w5882 , w12532 );
nor ( w5884 , w5883 , w5845 );
and ( w5885 , w5884 , w12037 );
not ( w5886 , w5885 );
and ( w5887 , w5886 , w5183 );
nor ( w5888 , w5887 , w2735 );
not ( w5889 , w5888 );
and ( w5890 , w5889 , w2582 );
not ( w5891 , w5890 );
and ( w5892 , w5891 , w2624 );
and ( w5893 , w5892 , w2587 );
nor ( w5894 , w5893 , w2575 );
and ( w5895 , w5894 , w6110 );
and ( w5896 , w255 , w5895 );
nor ( w5897 , w5896 , w5196 );
not ( w5898 , w2994 );
and ( w5899 , w5897 , w5898 );
and ( w5900 , w5899 , w20 );
and ( w5901 , w5900 , w11166 );
and ( w5902 , w20 , w5901 );
not ( w5903 , w5902 );
and ( w5904 , w5903 , w5105 );
and ( w5905 , w5904 , w5856 );
nor ( w5906 , w5905 , w310 );
nor ( w5907 , w5906 , w308 );
nor ( w5908 , w5907 , w5845 );
and ( w5909 , w5908 , w12037 );
not ( w5910 , w5909 );
and ( w5911 , w5910 , w5183 );
nor ( w5912 , w5911 , w2735 );
not ( w5913 , w5912 );
and ( w5914 , w5913 , w2582 );
not ( w5915 , w5914 );
and ( w5916 , w5915 , w2624 );
and ( w5917 , w5916 , w2587 );
nor ( w5918 , w5917 , w2575 );
and ( w5919 , w5918 , w6110 );
not ( w5920 , w5919 );
and ( w5921 , w5575 , w5920 );
and ( w5922 , w5921 , w12037 );
not ( w5923 , w5922 );
and ( w5924 , w5923 , w5183 );
nor ( w5925 , w5924 , w2735 );
not ( w5926 , w5925 );
and ( w5927 , w5926 , w2582 );
not ( w5928 , w5927 );
and ( w5929 , w5928 , w2587 );
nor ( w5930 , w5929 , w2575 );
and ( w5931 , w5930 , w6110 );
not ( w5932 , w5217 );
and ( w5933 , w5932 , w5931 );
and ( w5934 , w5933 , w12532 );
nor ( w5935 , w5934 , w5919 );
and ( w5936 , w5935 , w12037 );
not ( w5937 , w5936 );
and ( w5938 , w5937 , w5183 );
nor ( w5939 , w5938 , w2735 );
not ( w5940 , w5939 );
and ( w5941 , w5940 , w2582 );
not ( w5942 , w5941 );
and ( w5943 , w5942 , w2624 );
and ( w5944 , w5943 , w2587 );
nor ( w5945 , w5944 , w2575 );
and ( w5946 , w5945 , w6110 );
nor ( w5947 , w5213 , w5946 );
and ( w5948 , w5947 , w5968 );
and ( w5949 , w5948 , w2624 );
and ( w5950 , w5949 , w2587 );
nor ( w5951 , w5950 , w2575 );
nor ( w5952 , w5951 , w19 );
not ( w5953 , w5952 );
and ( w5954 , w5953 , w5678 );
not ( w5955 , w5954 );
and ( w5956 , w5955 , w308 );
and ( w5957 , w5956 , w310 );
and ( w5958 , w5957 , w11852 );
and ( w5959 , w5958 , w310 );
and ( w5960 , w5355 , w6008 );
nor ( w5961 , w5960 , w5946 );
and ( w5962 , w5961 , w5968 );
nor ( w5963 , w5962 , w2575 );
nor ( w5964 , w5963 , w48 );
nor ( w5965 , w5964 , w2592 );
and ( w5966 , w5965 , w12142 );
nor ( w5967 , w5966 , w5946 );
not ( w5968 , w2735 );
and ( w5969 , w5967 , w5968 );
and ( w5970 , w5969 , w2624 );
and ( w5971 , w5970 , w2587 );
nor ( w5972 , w5971 , w2575 );
and ( w5973 , w5972 , w6110 );
nor ( w5974 , w5973 , g31 );
nor ( w5975 , w5974 , g31 );
not ( w5976 , w5975 );
and ( w5977 , w5976 , w384 );
nor ( w5978 , w5966 , w255 );
nor ( w5979 , w5978 , w5578 );
not ( w5980 , w5979 );
and ( w5981 , w5980 , w308 );
and ( w5982 , w5981 , w11852 );
and ( w5983 , w5982 , w12717 );
not ( w5984 , w5946 );
and ( w5985 , w5983 , w5984 );
and ( w5986 , w5985 , w12037 );
not ( w5987 , w5986 );
and ( w5988 , w5987 , w5183 );
nor ( w5989 , w5988 , w2735 );
not ( w5990 , w5989 );
and ( w5991 , w5990 , w2582 );
not ( w5992 , w5991 );
and ( w5993 , w5992 , w2624 );
and ( w5994 , w5993 , w2587 );
nor ( w5995 , w5994 , w2575 );
and ( w5996 , w5995 , w6110 );
not ( w5997 , w5977 );
and ( w5998 , w5997 , w5996 );
and ( w5999 , w5998 , w8848 );
and ( w6000 , w5265 , w5189 );
and ( w6001 , w6000 , w5532 );
and ( w6002 , w6001 , w5183 );
not ( w6003 , w2575 );
and ( w6004 , w6002 , w6003 );
and ( w6005 , w2589 , w6004 );
and ( w6006 , w6005 , w19 );
and ( w6007 , w6006 , w2775 );
not ( w6008 , w5212 );
and ( w6009 , w6007 , w6008 );
nor ( w6010 , w6009 , w5946 );
nor ( w6011 , w6010 , w2592 );
and ( w6012 , w6011 , w5183 );
nor ( w6013 , w6012 , w2735 );
not ( w6014 , w6013 );
and ( w6015 , w6014 , w2582 );
not ( w6016 , w6015 );
and ( w6017 , w6016 , w2624 );
and ( w6018 , w6017 , w2587 );
nor ( w6019 , w6018 , w2575 );
and ( w6020 , w6019 , w6110 );
nor ( w6021 , w5999 , w6020 );
and ( w6022 , w6021 , w5365 );
and ( w6023 , w6022 , w12919 );
and ( w6024 , w12921 , w6023 );
not ( w6025 , w6024 );
and ( w6026 , w6025 , w2775 );
and ( w6027 , w6026 , w5532 );
nor ( w6028 , w6027 , w2961 );
and ( w6029 , w6028 , w12498 );
nor ( w6030 , w6029 , w5212 );
nor ( w6031 , w6030 , w5946 );
not ( w6032 , w6031 );
and ( w6033 , w6032 , w5183 );
nor ( w6034 , w6033 , w2735 );
not ( w6035 , w6034 );
and ( w6036 , w6035 , w2582 );
not ( w6037 , w6036 );
and ( w6038 , w6037 , w2624 );
and ( w6039 , w6038 , w2587 );
nor ( w6040 , w6039 , w2575 );
and ( w6041 , w6040 , w6110 );
not ( w6042 , w5959 );
and ( w6043 , w6042 , w6041 );
nor ( w6044 , w6043 , w18 );
and ( w6045 , w12921 , w6044 );
not ( w6046 , w6045 );
and ( w6047 , w6046 , w2775 );
and ( w6048 , w6047 , w5532 );
nor ( w6049 , w6048 , w377 );
nor ( w6050 , w6049 , w5212 );
nor ( w6051 , w6050 , w5946 );
and ( w6052 , w6051 , w12037 );
not ( w6053 , w6052 );
and ( w6054 , w6053 , w5183 );
nor ( w6055 , w6054 , w2735 );
not ( w6056 , w6055 );
and ( w6057 , w6056 , w2582 );
not ( w6058 , w6057 );
and ( w6059 , w6058 , w2624 );
and ( w6060 , w6059 , w2587 );
nor ( w6061 , w6060 , w2575 );
and ( w6062 , w6061 , w6110 );
nor ( w6063 , w5206 , w6062 );
not ( w6064 , w6063 );
and ( w6065 , w6064 , w5532 );
nor ( w6066 , w6065 , w312 );
not ( w6067 , w6066 );
and ( w6068 , w6067 , w5183 );
nor ( w6069 , w6068 , w2735 );
not ( w6070 , w6069 );
and ( w6071 , w6070 , w2582 );
not ( w6072 , w6071 );
and ( w6073 , w6072 , w2587 );
nor ( w6074 , w6073 , w2575 );
and ( w6075 , w6074 , w6110 );
and ( w6076 , w5202 , w6075 );
and ( w6077 , w6076 , w11166 );
nor ( w6078 , w6077 , w2961 );
nor ( w6079 , w6078 , w5212 );
nor ( w6080 , w6079 , w5946 );
not ( w6081 , w6080 );
and ( w6082 , w6081 , w5183 );
nor ( w6083 , w6082 , w2735 );
not ( w6084 , w6083 );
and ( w6085 , w6084 , w2582 );
not ( w6086 , w6085 );
and ( w6087 , w6086 , w2624 );
and ( w6088 , w6087 , w2587 );
nor ( w6089 , w6088 , w2575 );
and ( w6090 , w6089 , w6110 );
and ( w6091 , w19 , w6090 );
nor ( w6092 , w6091 , w2994 );
and ( w6093 , w20 , w6092 );
not ( w6094 , w6093 );
and ( w6095 , w6094 , w5105 );
and ( w6096 , w6095 , w6075 );
nor ( w6097 , w6096 , w2961 );
and ( w6098 , w6097 , w12498 );
nor ( w6099 , w6098 , w5212 );
nor ( w6100 , w6099 , w5946 );
not ( w6101 , w6100 );
and ( w6102 , w6101 , w5183 );
nor ( w6103 , w6102 , w2735 );
not ( w6104 , w6103 );
and ( w6105 , w6104 , w2582 );
not ( w6106 , w6105 );
and ( w6107 , w6106 , w2624 );
and ( w6108 , w6107 , w2587 );
nor ( w6109 , w6108 , w2575 );
not ( w6110 , w2592 );
and ( w6111 , w6109 , w6110 );
nor ( w6112 , w3169 , w212 );
not ( w6113 , w2586 );
and ( w6114 , w6112 , w6113 );
and ( w6115 , w6114 , w8 );
not ( w6116 , w6115 );
and ( w6117 , w6116 , w1 );
not ( w6118 , w6117 );
and ( w6119 , w6118 , w2643 );
nor ( w6120 , w3167 , w2586 );
not ( w6121 , w3169 );
and ( w6122 , w6120 , w6121 );
nor ( w6123 , w6122 , w2624 );
not ( w6124 , w6123 );
and ( w6125 , w6124 , w2587 );
and ( w6126 , w6119 , w6125 );
and ( w6127 , w6111 , w6130 );
and ( w6128 , w6148 , w6127 );
and ( w6129 , w6128 , w6111 );
not ( w6130 , w6126 );
and ( w6131 , w6129 , w6130 );
not ( w6132 , w6131 );
and ( w6133 , w6132 , w2587 );
nor ( w6134 , w2575 , w6133 );
and ( w6135 , w2664 , w7340 );
and ( w6136 , w6134 , w6135 );
nor ( w6137 , w10 , g3 );
not ( w6138 , g4 );
and ( w6139 , w6137 , w6138 );
nor ( w6140 , g5 , w8 );
and ( w6141 , w6140 , w12934 );
nor ( w6142 , w6141 , w66 );
nor ( w6143 , w11 , w6133 );
not ( w6144 , w8 );
and ( w6145 , w6143 , w6144 );
nor ( w6146 , w6145 , w2551 );
nor ( w6147 , w6146 , w6133 );
not ( w6148 , w14 );
and ( w6149 , w6147 , w6148 );
and ( w6150 , w6149 , w7340 );
and ( w6151 , w6142 , w6539 );
not ( w6152 , w6139 );
and ( w6153 , w6152 , w6151 );
and ( w6154 , w6153 , w6539 );
and ( w6155 , w1629 , w6539 );
and ( w6156 , w6155 , w12934 );
nor ( w6157 , w6156 , g5 );
and ( w6158 , w6157 , w12934 );
not ( w6159 , w6158 );
and ( w6160 , w6154 , w6159 );
and ( w6161 , w6160 , w11217 );
and ( w6162 , w6161 , w13211 );
not ( w6163 , w6162 );
and ( w6164 , w6163 , w6136 );
and ( w6165 , w6136 , w11217 );
not ( w6166 , w6165 );
and ( w6167 , w6166 , w6160 );
nor ( w6168 , w6167 , g33 );
and ( w6169 , w6136 , w7340 );
and ( w6170 , w7340 , g36 );
not ( w6171 , w6170 );
and ( w6172 , w6171 , w6160 );
not ( w6173 , w6172 );
and ( w6174 , w6173 , g11 );
and ( w6175 , w6160 , w13331 );
and ( w6176 , w6175 , w13333 );
nor ( w6177 , w6176 , w6133 );
and ( w6178 , w7340 , g39 );
and ( w6179 , w6178 , w6169 );
not ( w6180 , w6179 );
and ( w6181 , w6180 , w6160 );
not ( w6182 , w6181 );
and ( w6183 , w6182 , g13 );
nor ( w6184 , w6183 , w6174 );
and ( w6185 , w6798 , w6169 );
and ( w6186 , w6185 , w6136 );
and ( w6187 , w6134 , w13331 );
not ( w6188 , w6187 );
and ( w6189 , w6188 , w6160 );
nor ( w6190 , w6189 , g29 );
nor ( w6191 , w6186 , w6190 );
and ( w6192 , w6191 , w7354 );
and ( w6193 , w6136 , w6953 );
and ( w6194 , w6169 , w6135 );
and ( w6195 , w6194 , w6134 );
and ( w6196 , w6195 , w6136 );
not ( w6197 , g41 );
and ( w6198 , w6197 , w6160 );
and ( w6199 , w6205 , g15 );
not ( w6200 , w6199 );
and ( w6201 , w6200 , w6160 );
and ( w6202 , w6201 , w9053 );
not ( w6203 , w6202 );
and ( w6204 , w6203 , g17 );
not ( w6205 , w6198 );
and ( w6206 , w6205 , g40 );
and ( w6207 , w6206 , g15 );
not ( w6208 , w6207 );
and ( w6209 , w6208 , w6160 );
not ( w6210 , w6204 );
and ( w6211 , w6210 , w6209 );
not ( w6212 , w6211 );
and ( w6213 , w6196 , w6212 );
and ( w6214 , w6213 , w6134 );
and ( w6215 , w9195 , w6160 );
not ( w6216 , w6215 );
and ( w6217 , w6216 , g19 );
nor ( w6218 , w6214 , w6217 );
not ( w6219 , w6218 );
and ( w6220 , w6219 , w6136 );
not ( w6221 , w6217 );
and ( w6222 , w6221 , w6211 );
and ( w6223 , w6220 , w6695 );
and ( w6224 , w6223 , w6136 );
and ( w6225 , w6224 , w6134 );
and ( w6226 , w6225 , w6136 );
and ( w6227 , w6226 , w6134 );
and ( w6228 , w6227 , w6135 );
and ( w6229 , w6194 , w6136 );
and ( w6230 , w6229 , w6135 );
and ( w6231 , w6230 , w6134 );
and ( w6232 , w6231 , w6135 );
and ( w6233 , w6232 , w6134 );
and ( w6234 , w6134 , w6196 );
and ( w6235 , w6234 , w6136 );
and ( w6236 , w6235 , w6135 );
and ( w6237 , w6236 , w6134 );
and ( w6238 , w6233 , w6237 );
and ( w6239 , w6238 , w6134 );
and ( w6240 , w6239 , w6136 );
and ( w6241 , w6240 , w6134 );
and ( w6242 , w6241 , w6135 );
and ( w6243 , w6228 , w6242 );
and ( w6244 , w6160 , g37 );
and ( w6245 , w6244 , g19 );
not ( w6246 , w6245 );
and ( w6247 , w6246 , w6136 );
nor ( w6248 , w6133 , g40 );
not ( w6249 , w6248 );
and ( w6250 , w6249 , w6160 );
nor ( w6251 , w6250 , g17 );
and ( w6252 , w6169 , w6251 );
and ( w6253 , w6160 , g41 );
and ( w6254 , w6253 , g15 );
not ( w6255 , w6254 );
and ( w6256 , w6255 , w6134 );
and ( w6257 , w6136 , w6256 );
and ( w6258 , w6160 , g40 );
and ( w6259 , w6258 , g17 );
not ( w6260 , w6259 );
and ( w6261 , w6260 , w6134 );
and ( w6262 , w6261 , w6256 );
and ( w6263 , w6257 , w6262 );
nor ( w6264 , w6252 , w6263 );
not ( w6265 , w6264 );
and ( w6266 , w6247 , w6265 );
nor ( w6267 , w6243 , w6266 );
not ( w6268 , w6267 );
and ( w6269 , w6268 , w6136 );
and ( w6270 , w7340 , g42 );
not ( w6271 , w6270 );
and ( w6272 , w6271 , w6160 );
not ( w6273 , w6272 );
and ( w6274 , w6273 , g21 );
nor ( w6275 , w6269 , w6274 );
not ( w6276 , w6275 );
and ( w6277 , w6276 , w6136 );
and ( w6278 , w6277 , w6135 );
and ( w6279 , w6278 , w6134 );
and ( w6280 , w7340 , g43 );
not ( w6281 , w6280 );
and ( w6282 , w6281 , w6160 );
not ( w6283 , w6282 );
and ( w6284 , w6283 , g23 );
nor ( w6285 , w6279 , w6284 );
and ( w6286 , w6215 , w9197 );
not ( w6287 , w6286 );
and ( w6288 , w6287 , w6136 );
and ( w6289 , w6160 , w9053 );
and ( w6290 , w6289 , w9049 );
not ( w6291 , w6290 );
and ( w6292 , w6291 , g41 );
not ( w6293 , w6292 );
and ( w6294 , w6293 , w6160 );
not ( w6295 , w6294 );
and ( w6296 , w6295 , g15 );
nor ( w6297 , w6296 , w6217 );
not ( w6298 , w6289 );
and ( w6299 , w6298 , g17 );
not ( w6300 , w6299 );
and ( w6301 , w6297 , w6300 );
and ( w6302 , w6288 , w6640 );
and ( w6303 , w6302 , w6136 );
not ( w6304 , w6303 );
and ( w6305 , w6304 , w6160 );
and ( w6306 , w6305 , w9354 );
nor ( w6307 , w6306 , w6133 );
and ( w6308 , w6307 , g21 );
and ( w6309 , w6288 , g42 );
not ( w6310 , w6309 );
and ( w6311 , w6310 , w6160 );
nor ( w6312 , w6311 , w6301 );
and ( w6313 , w6312 , w6136 );
nor ( w6314 , w6308 , w6313 );
nor ( w6315 , w6285 , w6314 );
and ( w6316 , w6315 , w6136 );
and ( w6317 , w6316 , w6135 );
nor ( w6318 , w6317 , w6284 );
not ( w6319 , w6318 );
and ( w6320 , w6319 , w6169 );
and ( w6321 , w6320 , w6136 );
and ( w6322 , w6321 , w6135 );
and ( w6323 , w6160 , w9380 );
and ( w6324 , w6323 , w13321 );
nor ( w6325 , w6324 , w6133 );
and ( w6326 , w6322 , w6325 );
and ( w6327 , w6326 , w6136 );
and ( w6328 , w6160 , w12962 );
and ( w6329 , w6328 , w12964 );
not ( w6330 , w6329 );
and ( w6331 , w6330 , w6136 );
and ( w6332 , w6327 , w6331 );
and ( w6333 , w6332 , w6136 );
and ( w6334 , w7340 , g38 );
not ( w6335 , w6334 );
and ( w6336 , w6335 , w6160 );
not ( w6337 , w6336 );
and ( w6338 , w6337 , g25 );
nor ( w6339 , w6333 , w6338 );
not ( w6340 , w6339 );
and ( w6341 , w6340 , w6135 );
and ( w6342 , w6341 , w6136 );
and ( w6343 , w6136 , g44 );
not ( w6344 , w6343 );
and ( w6345 , w6344 , w6160 );
not ( w6346 , w6345 );
and ( w6347 , w6346 , g27 );
nor ( w6348 , w6342 , w6347 );
not ( w6349 , w6348 );
and ( w6350 , w6349 , w6169 );
and ( w6351 , w6350 , w6136 );
and ( w6352 , w6351 , w6135 );
and ( w6353 , w6352 , w6134 );
and ( w6354 , w6353 , w6136 );
and ( w6355 , w6354 , w6135 );
and ( w6356 , w6355 , w6134 );
and ( w6357 , w6356 , w6136 );
nor ( w6358 , w6133 , g42 );
and ( w6359 , w6358 , w9356 );
not ( w6360 , w6359 );
and ( w6361 , w6360 , w6160 );
and ( w6362 , w6361 , g37 );
and ( w6363 , w6362 , g19 );
not ( w6364 , w6363 );
and ( w6365 , w6364 , w6134 );
nor ( w6366 , w6133 , g37 );
not ( w6367 , w6366 );
and ( w6368 , w6367 , w6160 );
nor ( w6369 , w6368 , g19 );
nor ( w6370 , w6369 , w6251 );
not ( w6371 , w6370 );
and ( w6372 , w6371 , w6134 );
nor ( w6373 , w6372 , w6262 );
not ( w6374 , w6373 );
and ( w6375 , w6374 , w6134 );
and ( w6376 , w6375 , w7340 );
and ( w6377 , w6376 , w9354 );
not ( w6378 , w6377 );
and ( w6379 , w6378 , w6160 );
and ( w6380 , w6379 , g21 );
nor ( w6381 , w6369 , w6262 );
not ( w6382 , w6251 );
and ( w6383 , w6381 , w6382 );
and ( w6384 , w6383 , w6160 );
and ( w6385 , w6384 , g42 );
nor ( w6386 , w6385 , w6133 );
and ( w6387 , w6386 , w6134 );
not ( w6388 , w6380 );
and ( w6389 , w6388 , w6387 );
and ( w6390 , w6365 , w6389 );
and ( w6391 , w6390 , w6237 );
nor ( w6392 , w6133 , g43 );
and ( w6393 , w6392 , w13321 );
not ( w6394 , w6393 );
and ( w6395 , w6394 , w6160 );
not ( w6396 , w6391 );
and ( w6397 , w6396 , w6395 );
not ( w6398 , w6397 );
and ( w6399 , w6398 , w6134 );
and ( w6400 , w6990 , w6301 );
not ( w6401 , w6400 );
and ( w6402 , w6401 , w6136 );
and ( w6403 , w6402 , w6637 );
nor ( w6404 , w6403 , w6274 );
not ( w6405 , w6404 );
and ( w6406 , w6405 , w6136 );
and ( w6407 , w6406 , w6135 );
and ( w6408 , w6407 , w6237 );
and ( w6409 , w6408 , w6136 );
and ( w6410 , w6409 , w6134 );
nor ( w6411 , w6410 , w6284 );
not ( w6412 , w6411 );
and ( w6413 , w6412 , w6169 );
and ( w6414 , w6413 , w6136 );
and ( w6415 , w6160 , g44 );
not ( w6416 , w6415 );
and ( w6417 , w6416 , g44 );
nor ( w6418 , w6417 , w6150 );
and ( w6419 , w6418 , g27 );
not ( w6420 , w6419 );
and ( w6421 , w6420 , g27 );
and ( w6422 , g44 , w6539 );
and ( w6423 , w6422 , g27 );
not ( w6424 , w6423 );
and ( w6425 , w6424 , w6134 );
nor ( w6426 , w6421 , w6425 );
not ( w6427 , w6331 );
and ( w6428 , w6426 , w6427 );
not ( w6429 , w6428 );
and ( w6430 , w6429 , w6136 );
nor ( w6431 , w6430 , w6347 );
not ( w6432 , w6431 );
and ( w6433 , w6432 , w6136 );
and ( w6434 , w6433 , w6135 );
and ( w6435 , w6434 , w6134 );
and ( w6436 , w6435 , w6136 );
and ( w6437 , w6436 , w6135 );
and ( w6438 , w6437 , w6134 );
and ( w6439 , w6438 , w6136 );
and ( w6440 , w6160 , w8986 );
and ( w6441 , w6440 , w13050 );
not ( w6442 , w6441 );
and ( w6443 , w6442 , w6136 );
and ( w6444 , w6439 , w6443 );
and ( w6445 , w6134 , w8986 );
and ( w6446 , w6445 , w13050 );
not ( w6447 , w6446 );
and ( w6448 , w6447 , w6160 );
not ( w6449 , w6444 );
and ( w6450 , w6449 , w6448 );
not ( w6451 , w6450 );
and ( w6452 , w6451 , w6135 );
and ( w6453 , w6452 , w6134 );
and ( w6454 , w6414 , w6453 );
and ( w6455 , w6454 , w6136 );
and ( w6456 , w6455 , w6135 );
and ( w6457 , w6456 , w6134 );
and ( w6458 , w6457 , w6136 );
and ( w6459 , w6458 , w6135 );
and ( w6460 , w6459 , w6134 );
and ( w6461 , w6460 , w6136 );
and ( w6462 , w6461 , w6443 );
not ( w6463 , w6462 );
and ( w6464 , w6463 , w6448 );
not ( w6465 , w6464 );
and ( w6466 , w6465 , w6135 );
and ( w6467 , w6466 , w6134 );
and ( w6468 , w6357 , w6467 );
and ( w6469 , w6468 , w6443 );
and ( w6470 , w6160 , w9010 );
and ( w6471 , w6470 , w13590 );
not ( w6472 , w6471 );
and ( w6473 , w6472 , w6136 );
and ( w6474 , w6469 , w6473 );
and ( w6475 , w6338 , w6134 );
nor ( w6476 , w6475 , w6347 );
not ( w6477 , w6476 );
and ( w6478 , w6477 , w6134 );
and ( w6479 , w6478 , w6136 );
and ( w6480 , w6136 , w6695 );
and ( w6481 , w6480 , w6134 );
nor ( w6482 , w6481 , w6274 );
not ( w6483 , w6482 );
and ( w6484 , w6483 , w6134 );
and ( w6485 , w6484 , w6136 );
nor ( w6486 , w6485 , w6284 );
not ( w6487 , w6486 );
and ( w6488 , w6487 , w6134 );
and ( w6489 , w6488 , w6136 );
and ( w6490 , w6489 , w6135 );
and ( w6491 , w6490 , w6136 );
and ( w6492 , w6491 , w6134 );
and ( w6493 , w6492 , w6136 );
nor ( w6494 , w6479 , w6493 );
and ( w6495 , w6160 , g43 );
and ( w6496 , w6495 , g23 );
nor ( w6497 , w6496 , w6133 );
not ( w6498 , w6497 );
and ( w6499 , w6498 , w6395 );
not ( w6500 , w6499 );
and ( w6501 , w6500 , w6134 );
and ( w6502 , w6501 , w6169 );
and ( w6503 , w6389 , w6135 );
and ( w6504 , w6503 , w6134 );
and ( w6505 , w6504 , w6135 );
and ( w6506 , w6505 , w6136 );
and ( w6507 , w6136 , w9195 );
not ( w6508 , w6507 );
and ( w6509 , w6508 , w6160 );
nor ( w6510 , w6509 , g19 );
and ( w6511 , w6136 , w9354 );
and ( w6512 , w6511 , w9356 );
not ( w6513 , w6512 );
and ( w6514 , w6513 , w6160 );
not ( w6515 , w6510 );
and ( w6516 , w6515 , w6514 );
not ( w6517 , w6266 );
and ( w6518 , w6516 , w6517 );
not ( w6519 , w6518 );
and ( w6520 , w6506 , w6519 );
not ( w6521 , w6520 );
and ( w6522 , w6521 , w6395 );
not ( w6523 , w6522 );
and ( w6524 , w6523 , w6169 );
and ( w6525 , w6524 , w6134 );
and ( w6526 , w6525 , w6136 );
and ( w6527 , w6502 , w6526 );
and ( w6528 , w6527 , w6136 );
and ( w6529 , w6528 , w6135 );
and ( w6530 , w6529 , w6134 );
and ( w6531 , w6136 , w12962 );
and ( w6532 , w6531 , w12964 );
not ( w6533 , w6532 );
and ( w6534 , w6533 , w6160 );
not ( w6535 , w6530 );
and ( w6536 , w6535 , w6534 );
not ( w6537 , w6536 );
and ( w6538 , w6537 , w6134 );
not ( w6539 , w6150 );
and ( w6540 , g38 , w6539 );
and ( w6541 , w6540 , g25 );
not ( w6542 , w6541 );
and ( w6543 , w6542 , w6134 );
and ( w6544 , w6538 , w6543 );
and ( w6545 , w6160 , g38 );
not ( w6546 , w6545 );
and ( w6547 , w6546 , g38 );
nor ( w6548 , w6547 , w6150 );
and ( w6549 , w6548 , g25 );
not ( w6550 , w6549 );
and ( w6551 , w6550 , g25 );
nor ( w6552 , w6544 , w6551 );
not ( w6553 , w6552 );
and ( w6554 , w6553 , w6134 );
and ( w6555 , w6554 , w6136 );
and ( w6556 , w6555 , w6425 );
nor ( w6557 , w6556 , w6421 );
and ( w6558 , w6494 , w6557 );
and ( w6559 , w6558 , w6448 );
and ( w6560 , w6347 , w6960 );
and ( w6561 , w6169 , w6284 );
and ( w6562 , w6960 , w6136 );
and ( w6563 , w6562 , w6473 );
not ( w6564 , w6314 );
and ( w6565 , w6134 , w6564 );
and ( w6566 , w6565 , w6136 );
and ( w6567 , w6566 , w6169 );
and ( w6568 , w6567 , w6325 );
nor ( w6569 , w6568 , w6338 );
not ( w6570 , w6569 );
and ( w6571 , w6570 , w6169 );
and ( w6572 , w6571 , w6473 );
and ( w6573 , w6331 , w6572 );
and ( w6574 , w6563 , w6573 );
and ( w6575 , w6574 , w6443 );
not ( w6576 , w6575 );
and ( w6577 , w6576 , w6448 );
not ( w6578 , w6577 );
and ( w6579 , w6578 , w6136 );
and ( w6580 , w6579 , w6135 );
and ( w6581 , w6580 , w6134 );
and ( w6582 , w6581 , w6960 );
and ( w6583 , w6582 , w6134 );
and ( w6584 , w6583 , w6136 );
and ( w6585 , w6584 , w6134 );
and ( w6586 , w6585 , w6497 );
and ( w6587 , w6586 , w6331 );
and ( w6588 , w6587 , w6136 );
and ( w6589 , w6588 , w6443 );
and ( w6590 , w6589 , w6473 );
and ( w6591 , w6590 , w6136 );
and ( w6592 , w6591 , w6135 );
and ( w6593 , w6592 , w6134 );
nor ( w6594 , w6561 , w6593 );
nor ( w6595 , w6594 , w6559 );
and ( w6596 , w6595 , w6331 );
and ( w6597 , w6596 , w6136 );
and ( w6598 , w6597 , w6443 );
and ( w6599 , w6598 , w6473 );
nor ( w6600 , w6560 , w6599 );
not ( w6601 , w6600 );
and ( w6602 , w6601 , w6136 );
and ( w6603 , w6602 , w6443 );
and ( w6604 , w6603 , w6473 );
and ( w6605 , w6474 , w6604 );
and ( w6606 , w6169 , w6134 );
and ( w6607 , w6606 , w7340 );
and ( w6608 , w6607 , w6134 );
and ( w6609 , w6562 , w6608 );
and ( w6610 , w6609 , w6134 );
and ( w6611 , w6610 , w6136 );
and ( w6612 , w6611 , w7340 );
and ( w6613 , w6612 , w6134 );
and ( w6614 , w6613 , w6174 );
nor ( w6615 , w6614 , w6183 );
not ( w6616 , w6615 );
and ( w6617 , w6616 , w6134 );
nor ( w6618 , w6617 , w6177 );
not ( w6619 , w6618 );
and ( w6620 , w6619 , w6134 );
and ( w6621 , w6620 , w6136 );
and ( w6622 , w6621 , w7340 );
and ( w6623 , w6622 , w6134 );
and ( w6624 , w6623 , w6953 );
and ( w6625 , w6134 , g48 );
not ( w6626 , w6625 );
and ( w6627 , w6626 , w6160 );
not ( w6628 , w6627 );
and ( w6629 , w6628 , g31 );
and ( w6630 , w6624 , w6629 );
and ( w6631 , w6606 , w6136 );
and ( w6632 , w6631 , w6467 );
and ( w6633 , w6632 , w6443 );
and ( w6634 , w6633 , w6473 );
and ( w6635 , w6634 , w6347 );
and ( w6636 , w6169 , w6284 );
not ( w6637 , w6285 );
and ( w6638 , w6637 , w6136 );
and ( w6639 , w6638 , w6135 );
not ( w6640 , w6301 );
and ( w6641 , w6639 , w6640 );
and ( w6642 , w6641 , w6136 );
and ( w6643 , w6642 , w6135 );
and ( w6644 , w6643 , w6169 );
and ( w6645 , w6644 , w6325 );
nor ( w6646 , w6645 , w6338 );
not ( w6647 , w6646 );
and ( w6648 , w6647 , w6134 );
and ( w6649 , w6237 , w6136 );
and ( w6650 , w6649 , w6135 );
and ( w6651 , w6648 , w6650 );
and ( w6652 , w6651 , w6134 );
and ( w6653 , w6652 , w6136 );
and ( w6654 , w6653 , w6134 );
and ( w6655 , w6654 , w6497 );
and ( w6656 , w6655 , w6135 );
nor ( w6657 , w6656 , w6274 );
not ( w6658 , w6657 );
and ( w6659 , w6658 , w6136 );
and ( w6660 , w6659 , w6135 );
and ( w6661 , w6660 , w6650 );
and ( w6662 , w6661 , w6134 );
and ( w6663 , w6662 , w6497 );
and ( w6664 , w6663 , w6135 );
nor ( w6665 , w6636 , w6664 );
not ( w6666 , w6665 );
and ( w6667 , w6666 , w6135 );
and ( w6668 , w6667 , w6325 );
nor ( w6669 , w6668 , w6338 );
not ( w6670 , w6669 );
and ( w6671 , w6670 , w6136 );
and ( w6672 , w6671 , w6169 );
and ( w6673 , w6672 , w6136 );
and ( w6674 , w6673 , w6135 );
and ( w6675 , w6674 , w6134 );
and ( w6676 , w6675 , w7340 );
and ( w6677 , w6676 , w6134 );
and ( w6678 , w6677 , w6136 );
and ( w6679 , w6678 , w6467 );
and ( w6680 , w6679 , w6331 );
and ( w6681 , w6680 , w6599 );
and ( w6682 , w6681 , w6135 );
and ( w6683 , w6682 , w6136 );
and ( w6684 , w6683 , w6443 );
and ( w6685 , w6684 , w6473 );
and ( w6686 , w6685 , w6135 );
and ( w6687 , w6686 , w6134 );
and ( w6688 , w6687 , w6136 );
and ( w6689 , w6688 , w6135 );
and ( w6690 , w6136 , w6242 );
and ( w6691 , w6690 , w6134 );
and ( w6692 , w6691 , w6136 );
and ( w6693 , w6692 , w6228 );
and ( w6694 , w6693 , w6136 );
not ( w6695 , w6222 );
and ( w6696 , w6694 , w6695 );
and ( w6697 , w6696 , w6136 );
and ( w6698 , w6697 , w6134 );
and ( w6699 , w6698 , w6136 );
and ( w6700 , w6699 , w6134 );
nor ( w6701 , w6700 , w6284 );
not ( w6702 , w6701 );
and ( w6703 , w6702 , w6135 );
nor ( w6704 , w6703 , w6274 );
not ( w6705 , w6704 );
and ( w6706 , w6705 , w6135 );
and ( w6707 , w6706 , w6136 );
and ( w6708 , w6707 , w6135 );
and ( w6709 , w6708 , w6136 );
and ( w6710 , w6709 , w6169 );
and ( w6711 , w6710 , w6136 );
nor ( w6712 , w6711 , w6347 );
not ( w6713 , w6712 );
and ( w6714 , w6713 , w6136 );
nor ( w6715 , w6714 , w6338 );
not ( w6716 , w6715 );
and ( w6717 , w6716 , w6135 );
and ( w6718 , w6717 , w6169 );
and ( w6719 , w6718 , w6136 );
and ( w6720 , w6719 , w6135 );
and ( w6721 , w6720 , w6134 );
and ( w6722 , w6721 , w6135 );
and ( w6723 , w6722 , w6136 );
and ( w6724 , w6723 , w7340 );
and ( w6725 , w6724 , w6134 );
and ( w6726 , w6725 , w6136 );
and ( w6727 , w6726 , w6960 );
and ( w6728 , w6727 , w6136 );
not ( w6729 , w6728 );
and ( w6730 , w6729 , w6557 );
and ( w6731 , w6730 , w6448 );
not ( w6732 , w6731 );
and ( w6733 , w6732 , w6136 );
nor ( w6734 , w6572 , w6183 );
not ( w6735 , w6734 );
and ( w6736 , w6735 , w6134 );
and ( w6737 , w6736 , w6136 );
and ( w6738 , w6737 , w6134 );
and ( w6739 , w6738 , w6497 );
nor ( w6740 , w6739 , w6347 );
not ( w6741 , w6740 );
and ( w6742 , w6741 , w6443 );
nor ( w6743 , w6742 , w6183 );
not ( w6744 , w6743 );
and ( w6745 , w6744 , w6473 );
nor ( w6746 , w6745 , w6183 );
not ( w6747 , w6561 );
and ( w6748 , w6747 , w6746 );
not ( w6749 , w6748 );
and ( w6750 , w6749 , w6331 );
nor ( w6751 , w6750 , w6347 );
not ( w6752 , w6751 );
and ( w6753 , w6752 , w6443 );
nor ( w6754 , w6753 , w6183 );
not ( w6755 , w6754 );
and ( w6756 , w6755 , w6473 );
nor ( w6757 , w6756 , w6183 );
and ( w6758 , w6757 , w7356 );
not ( w6759 , w6758 );
and ( w6760 , w6759 , w6169 );
and ( w6761 , w6160 , g45 );
and ( w6762 , w6761 , g29 );
nor ( w6763 , w6762 , w6133 );
nor ( w6764 , w6760 , w6763 );
not ( w6765 , w6190 );
and ( w6766 , w6764 , w6765 );
nor ( w6767 , w6766 , w6133 );
and ( w6768 , w6767 , w6134 );
and ( w6769 , w6768 , w6135 );
and ( w6770 , w6769 , w6134 );
and ( w6771 , w6770 , w6136 );
nor ( w6772 , w6771 , w6183 );
not ( w6773 , w6772 );
and ( w6774 , w6733 , w6773 );
and ( w6775 , w6774 , w6136 );
nor ( w6776 , w6133 , g39 );
not ( w6777 , w6776 );
and ( w6778 , w6777 , w6160 );
nor ( w6779 , w6778 , g13 );
nor ( w6780 , w6775 , w6779 );
and ( w6781 , w6134 , g46 );
not ( w6782 , w6781 );
and ( w6783 , w6782 , w6160 );
not ( w6784 , w6783 );
and ( w6785 , w6784 , g9 );
and ( w6786 , w6780 , w7215 );
not ( w6787 , w6786 );
and ( w6788 , w6787 , w6135 );
and ( w6789 , w6788 , w6136 );
and ( w6790 , w6789 , w6135 );
and ( w6791 , w6790 , w6134 );
and ( w6792 , w6689 , w6791 );
and ( w6793 , w6792 , w6135 );
and ( w6794 , w6793 , w6134 );
nor ( w6795 , w6635 , w6794 );
not ( w6796 , w6795 );
and ( w6797 , w6796 , w6604 );
not ( w6798 , w6184 );
and ( w6799 , w6798 , w6608 );
and ( w6800 , w6799 , w6134 );
nor ( w6801 , w6800 , w6347 );
not ( w6802 , w6801 );
and ( w6803 , w6802 , w6136 );
and ( w6804 , w6803 , w6134 );
and ( w6805 , w6804 , w6136 );
nor ( w6806 , w6805 , w6443 );
not ( w6807 , w6806 );
and ( w6808 , w6807 , w6136 );
and ( w6809 , w6808 , w6134 );
and ( w6810 , w6134 , w6650 );
and ( w6811 , w6810 , w6135 );
and ( w6812 , w6811 , w6136 );
and ( w6813 , w6812 , w6543 );
nor ( w6814 , w6813 , w6551 );
not ( w6815 , w6814 );
and ( w6816 , w6815 , w6425 );
nor ( w6817 , w6816 , w6421 );
and ( w6818 , w6136 , w9010 );
and ( w6819 , w6818 , w13590 );
not ( w6820 , w6819 );
and ( w6821 , w6820 , w6160 );
and ( w6822 , w6817 , w6821 );
not ( w6823 , w6822 );
and ( w6824 , w6823 , w6135 );
and ( w6825 , w6824 , w6136 );
and ( w6826 , w6825 , w6134 );
and ( w6827 , w6826 , w6136 );
and ( w6828 , w6827 , w6134 );
and ( w6829 , w6828 , w7340 );
and ( w6830 , w6829 , w6134 );
and ( w6831 , w6830 , w6174 );
nor ( w6832 , w6831 , w6183 );
not ( w6833 , w6832 );
and ( w6834 , w6833 , w6134 );
and ( w6835 , w6834 , w7340 );
and ( w6836 , w6835 , w6134 );
and ( w6837 , w6836 , w6190 );
and ( w6838 , w6284 , w6134 );
and ( w6839 , w6838 , w6136 );
and ( w6840 , w6839 , w6331 );
nor ( w6841 , w6840 , w6338 );
not ( w6842 , w6841 );
and ( w6843 , w6842 , w6134 );
and ( w6844 , w6843 , w6136 );
and ( w6845 , w6844 , w6473 );
nor ( w6846 , w6845 , w6183 );
and ( w6847 , w6846 , w7356 );
not ( w6848 , w6847 );
and ( w6849 , w6848 , w6169 );
and ( w6850 , w6849 , w6467 );
and ( w6851 , w6850 , w6136 );
and ( w6852 , w6851 , w7340 );
and ( w6853 , w6852 , w6134 );
and ( w6854 , w6853 , w6177 );
not ( w6855 , w6176 );
and ( w6856 , w6855 , w6136 );
and ( w6857 , w6856 , w6169 );
and ( w6858 , w6857 , w6174 );
nor ( w6859 , w6183 , w6338 );
not ( w6860 , w6859 );
and ( w6861 , w6860 , w6134 );
and ( w6862 , w6861 , w6136 );
and ( w6863 , w6862 , w6473 );
nor ( w6864 , w6863 , w6183 );
and ( w6865 , w6864 , w6448 );
and ( w6866 , w6865 , w7354 );
not ( w6867 , w6858 );
and ( w6868 , w6867 , w6866 );
not ( w6869 , w6868 );
and ( w6870 , w6467 , w6869 );
and ( w6871 , w6870 , w7340 );
and ( w6872 , w6871 , w6134 );
and ( w6873 , w6872 , w6177 );
and ( w6874 , w7340 , g45 );
not ( w6875 , w6874 );
and ( w6876 , w6875 , w6160 );
not ( w6877 , w6876 );
and ( w6878 , w6877 , g29 );
nor ( w6879 , w6873 , w6878 );
not ( w6880 , w6879 );
and ( w6881 , w6880 , w6135 );
and ( w6882 , w6881 , w6134 );
and ( w6883 , w6882 , w6136 );
nor ( w6884 , w6883 , w6779 );
and ( w6885 , w6884 , w7215 );
not ( w6886 , w6885 );
and ( w6887 , w6886 , w6135 );
and ( w6888 , w6887 , w6791 );
and ( w6889 , w6888 , w6136 );
and ( w6890 , w6889 , w6135 );
and ( w6891 , w6890 , w6134 );
and ( w6892 , w6443 , w6891 );
nor ( w6893 , w6892 , w6183 );
and ( w6894 , w6893 , w7356 );
not ( w6895 , w6894 );
and ( w6896 , w6895 , w6169 );
and ( w6897 , w6896 , w6136 );
and ( w6898 , w6897 , w7340 );
and ( w6899 , w6898 , w6134 );
and ( w6900 , w6899 , w6177 );
nor ( w6901 , w6900 , w6878 );
not ( w6902 , w6901 );
and ( w6903 , w6902 , w6135 );
and ( w6904 , w6903 , w6134 );
and ( w6905 , w6904 , w6136 );
nor ( w6906 , w6905 , w6779 );
and ( w6907 , w6906 , w7215 );
not ( w6908 , w6907 );
and ( w6909 , w6908 , w6135 );
and ( w6910 , w6909 , w6791 );
and ( w6911 , w6910 , w6136 );
and ( w6912 , w6911 , w6135 );
and ( w6913 , w6912 , w6134 );
nor ( w6914 , w6854 , w6913 );
and ( w6915 , w6467 , w6604 );
nor ( w6916 , w6915 , w6913 );
nor ( w6917 , w6916 , w6133 );
and ( w6918 , w6917 , w6134 );
and ( w6919 , w6918 , w6177 );
and ( w6920 , w6356 , w6467 );
and ( w6921 , w6920 , w6604 );
and ( w6922 , w6921 , w6136 );
and ( w6923 , w6922 , w6443 );
and ( w6924 , w6923 , w6473 );
and ( w6925 , w6136 , g33 );
nor ( w6926 , w6925 , w6168 );
not ( w6927 , w6926 );
and ( w6928 , w6927 , w6134 );
and ( w6929 , w6928 , w6136 );
and ( w6930 , w6562 , w6929 );
and ( w6931 , w6930 , w6134 );
and ( w6932 , w6931 , w6136 );
and ( w6933 , w6932 , w6134 );
and ( w6934 , w6933 , w6136 );
and ( w6935 , w6934 , w6791 );
and ( w6936 , w6935 , w6136 );
and ( w6937 , w6929 , w6936 );
and ( w6938 , w6937 , w6134 );
and ( w6939 , w6938 , w6136 );
and ( w6940 , w6939 , w6134 );
and ( w6941 , w6940 , w6169 );
and ( w6942 , w6941 , w7340 );
and ( w6943 , w6942 , w6134 );
and ( w6944 , w6943 , w6174 );
nor ( w6945 , w6944 , w6183 );
and ( w6946 , w6945 , w6160 );
and ( w6947 , w6946 , w13331 );
and ( w6948 , w6947 , w13333 );
nor ( w6949 , w6948 , w6133 );
and ( w6950 , w6949 , w6136 );
and ( w6951 , w6950 , w7340 );
and ( w6952 , w6951 , w6134 );
not ( w6953 , w6192 );
and ( w6954 , w6952 , w6953 );
and ( w6955 , w6954 , w6136 );
and ( w6956 , w6955 , w6134 );
and ( w6957 , w6956 , w6629 );
and ( w6958 , w6606 , w6467 );
and ( w6959 , w6958 , w6135 );
not ( w6960 , w6559 );
and ( w6961 , w6959 , w6960 );
and ( w6962 , w6961 , w6136 );
and ( w6963 , w6962 , w6347 );
nor ( w6964 , w6963 , w6794 );
not ( w6965 , w6964 );
and ( w6966 , w6965 , w6135 );
and ( w6967 , w6160 , g48 );
and ( w6968 , w6967 , g31 );
nor ( w6969 , w6968 , w6133 );
and ( w6970 , w6966 , w6969 );
and ( w6971 , w6970 , w6136 );
and ( w6972 , w6971 , w6443 );
and ( w6973 , w6972 , w6473 );
and ( w6974 , w6606 , w6174 );
nor ( w6975 , w6974 , w6183 );
not ( w6976 , w6975 );
and ( w6977 , w6976 , w6134 );
and ( w6978 , w6977 , w6136 );
and ( w6979 , w6978 , w6134 );
and ( w6980 , w6979 , w6136 );
not ( w6981 , w6821 );
and ( w6982 , w6980 , w6981 );
and ( w6983 , w6631 , w6174 );
nor ( w6984 , w6983 , w6183 );
not ( w6985 , w6984 );
and ( w6986 , w6985 , w6134 );
not ( w6987 , w6448 );
and ( w6988 , w6986 , w6987 );
and ( w6989 , w6274 , w6134 );
not ( w6990 , w6399 );
and ( w6991 , w6990 , w6395 );
and ( w6992 , w6991 , w6534 );
not ( w6993 , w6992 );
and ( w6994 , w6993 , w6237 );
and ( w6995 , w6994 , w6136 );
and ( w6996 , w6995 , w6543 );
nor ( w6997 , w6996 , w6551 );
not ( w6998 , w6997 );
and ( w6999 , w6998 , w6425 );
nor ( w7000 , w6999 , w6421 );
and ( w7001 , w7000 , w6821 );
not ( w7002 , w7001 );
and ( w7003 , w7002 , w6136 );
and ( w7004 , w7003 , w6134 );
and ( w7005 , w6399 , w6497 );
not ( w7006 , w7005 );
and ( w7007 , w7006 , w6534 );
and ( w7008 , w7007 , w6395 );
not ( w7009 , w7008 );
and ( w7010 , w7009 , w6134 );
and ( w7011 , w7010 , w6543 );
nor ( w7012 , w7011 , w6551 );
and ( w7013 , w7012 , w6448 );
not ( w7014 , w7013 );
and ( w7015 , w7014 , w6136 );
and ( w7016 , w7015 , w6425 );
nor ( w7017 , w7016 , w6421 );
and ( w7018 , w7017 , g9 );
not ( w7019 , w7018 );
and ( w7020 , w7019 , w6134 );
and ( w7021 , w7020 , w6136 );
and ( w7022 , w7021 , w6134 );
nor ( w7023 , w7022 , w6779 );
not ( w7024 , w7023 );
and ( w7025 , w7024 , w6136 );
and ( w7026 , w7025 , w6134 );
and ( w7027 , w7026 , w6135 );
and ( w7028 , w7027 , w6136 );
and ( w7029 , w7028 , w6135 );
and ( w7030 , w7029 , w6134 );
and ( w7031 , w7004 , w7030 );
and ( w7032 , w7031 , w6134 );
and ( w7033 , w7032 , w6136 );
and ( w7034 , w7033 , w6134 );
nor ( w7035 , w7034 , w6779 );
not ( w7036 , w7035 );
and ( w7037 , w7036 , w6135 );
and ( w7038 , w7037 , w6134 );
nor ( w7039 , w6989 , w7038 );
not ( w7040 , w6284 );
and ( w7041 , w7039 , w7040 );
not ( w7042 , w7041 );
and ( w7043 , w7042 , w6136 );
and ( w7044 , w7043 , w6169 );
and ( w7045 , w7044 , w6134 );
and ( w7046 , w7045 , w6136 );
and ( w7047 , w7046 , w6543 );
nor ( w7048 , w7047 , w6551 );
not ( w7049 , w7048 );
and ( w7050 , w7049 , w6425 );
not ( w7051 , w6557 );
and ( w7052 , w7050 , w7051 );
nor ( w7053 , w7052 , w6421 );
and ( w7054 , w7053 , w6821 );
not ( w7055 , w7054 );
and ( w7056 , w7055 , w6136 );
and ( w7057 , w7056 , w6134 );
and ( w7058 , w7057 , w6136 );
and ( w7059 , w7058 , w6134 );
and ( w7060 , w7059 , w6136 );
and ( w7061 , w7060 , w6134 );
and ( w7062 , w7061 , w6169 );
and ( w7063 , w7062 , w7340 );
and ( w7064 , w7063 , w6134 );
and ( w7065 , w7064 , w6174 );
and ( w7066 , w6561 , w6331 );
nor ( w7067 , w7066 , w6183 );
not ( w7068 , w6338 );
and ( w7069 , w7067 , w7068 );
not ( w7070 , w7069 );
and ( w7071 , w7070 , w6134 );
and ( w7072 , w7071 , w6543 );
nor ( w7073 , w7072 , w6551 );
nor ( w7074 , w7073 , w6557 );
nor ( w7075 , w7074 , w6183 );
not ( w7076 , w7075 );
and ( w7077 , w7076 , w6443 );
nor ( w7078 , w7077 , w6183 );
not ( w7079 , w7065 );
and ( w7080 , w7079 , w7078 );
not ( w7081 , w7080 );
and ( w7082 , w7081 , w6443 );
not ( w7083 , w6968 );
and ( w7084 , w7083 , w6134 );
and ( w7085 , w7082 , w7084 );
nor ( w7086 , w7085 , w6878 );
not ( w7087 , w7086 );
and ( w7088 , w7087 , w6135 );
and ( w7089 , w7088 , w6134 );
and ( w7090 , w7089 , w6136 );
nor ( w7091 , w7090 , w6779 );
and ( w7092 , w7091 , w7215 );
not ( w7093 , w7092 );
and ( w7094 , w7093 , w6134 );
and ( w7095 , w7094 , w6135 );
and ( w7096 , w7095 , w6791 );
and ( w7097 , w7096 , w6136 );
and ( w7098 , w7097 , w6135 );
and ( w7099 , w7098 , w6134 );
nor ( w7100 , w6988 , w7099 );
not ( w7101 , w7100 );
and ( w7102 , w7101 , w7084 );
nor ( w7103 , w7102 , w6878 );
not ( w7104 , w7103 );
and ( w7105 , w7104 , w6135 );
and ( w7106 , w7105 , w6134 );
and ( w7107 , w7106 , w6136 );
nor ( w7108 , w7107 , w6785 );
not ( w7109 , w7108 );
and ( w7110 , w7109 , w6134 );
and ( w7111 , w7110 , w6791 );
and ( w7112 , w7111 , w6136 );
nor ( w7113 , w6982 , w7112 );
not ( w7114 , w7113 );
and ( w7115 , w7114 , w7084 );
nor ( w7116 , w7115 , w6878 );
not ( w7117 , w7116 );
and ( w7118 , w7117 , w6135 );
and ( w7119 , w7118 , w6134 );
and ( w7120 , w7119 , w6136 );
nor ( w7121 , w7120 , w6779 );
and ( w7122 , w7121 , w7215 );
not ( w7123 , w7122 );
and ( w7124 , w7123 , w6134 );
and ( w7125 , w7124 , w6135 );
and ( w7126 , w7125 , w6791 );
and ( w7127 , w7126 , w6136 );
and ( w7128 , w7127 , w6135 );
and ( w7129 , w7128 , w6134 );
nor ( w7130 , w6973 , w7129 );
not ( w7131 , w7130 );
and ( w7132 , w7131 , w6135 );
and ( w7133 , w7132 , w6134 );
and ( w7134 , w7133 , w6136 );
nor ( w7135 , w7134 , w6183 );
and ( w7136 , w7135 , w7215 );
not ( w7137 , w7136 );
and ( w7138 , w7137 , w6135 );
and ( w7139 , w7138 , w6791 );
and ( w7140 , w7139 , w6136 );
and ( w7141 , w7140 , w6135 );
and ( w7142 , w7141 , w6134 );
nor ( w7143 , w6957 , w7142 );
and ( w7144 , w7143 , w7263 );
not ( w7145 , w7144 );
and ( w7146 , w7145 , w6135 );
and ( w7147 , w7146 , w6134 );
and ( w7148 , w7147 , w6136 );
nor ( w7149 , w7148 , w6183 );
not ( w7150 , w7149 );
and ( w7151 , w7150 , w6136 );
nor ( w7152 , w7151 , w6785 );
not ( w7153 , w7152 );
and ( w7154 , w7153 , w6791 );
and ( w7155 , w7154 , w6136 );
nor ( w7156 , w6924 , w7155 );
not ( w7157 , w7156 );
and ( w7158 , w7157 , w6136 );
and ( w7159 , w7158 , w6629 );
nor ( w7160 , w7159 , w7142 );
and ( w7161 , w7160 , w7263 );
not ( w7162 , w7161 );
and ( w7163 , w7162 , w6135 );
and ( w7164 , w7163 , w6134 );
and ( w7165 , w7164 , w6136 );
and ( w7166 , w7165 , w6791 );
and ( w7167 , w7166 , w6135 );
and ( w7168 , w7167 , w6134 );
nor ( w7169 , w6919 , w7168 );
and ( w7170 , w7169 , w7263 );
not ( w7171 , w7170 );
and ( w7172 , w7171 , w6135 );
and ( w7173 , w7172 , w6134 );
and ( w7174 , w7173 , w6136 );
and ( w7175 , w7174 , w6791 );
not ( w7176 , w7175 );
and ( w7177 , w6914 , w7176 );
and ( w7178 , w7177 , w7263 );
not ( w7179 , w7178 );
and ( w7180 , w7179 , w6135 );
and ( w7181 , w7180 , w6134 );
and ( w7182 , w7181 , w6136 );
nor ( w7183 , w7182 , w6183 );
not ( w7184 , w6779 );
and ( w7185 , w7183 , w7184 );
and ( w7186 , w7185 , w7215 );
not ( w7187 , w7186 );
and ( w7188 , w7187 , w6135 );
and ( w7189 , w7188 , w6791 );
and ( w7190 , w7189 , w6136 );
and ( w7191 , w7190 , w6135 );
and ( w7192 , w7191 , w6134 );
nor ( w7193 , w6837 , w7192 );
not ( w7194 , w7193 );
and ( w7195 , w7194 , w6135 );
and ( w7196 , w7195 , w6136 );
and ( w7197 , w7196 , w6443 );
not ( w7198 , w7197 );
and ( w7199 , w7198 , w6448 );
not ( w7200 , w6913 );
and ( w7201 , w7199 , w7200 );
not ( w7202 , w7201 );
and ( w7203 , w7202 , w6969 );
and ( w7204 , w7203 , w7084 );
nor ( w7205 , w7204 , w7175 );
and ( w7206 , w7205 , w7263 );
not ( w7207 , w7206 );
and ( w7208 , w7207 , w6135 );
and ( w7209 , w7208 , w6134 );
and ( w7210 , w7209 , w6136 );
nor ( w7211 , w7210 , w6183 );
not ( w7212 , w7211 );
and ( w7213 , w7212 , w6136 );
nor ( w7214 , w7213 , w6779 );
not ( w7215 , w6785 );
and ( w7216 , w7214 , w7215 );
not ( w7217 , w7216 );
and ( w7218 , w7217 , w6134 );
and ( w7219 , w7218 , w6135 );
and ( w7220 , w7219 , w6791 );
and ( w7221 , w7220 , w6136 );
and ( w7222 , w7221 , w6135 );
and ( w7223 , w7222 , w6134 );
and ( w7224 , w6809 , w7223 );
nor ( w7225 , w7224 , w6913 );
not ( w7226 , w7225 );
and ( w7227 , w7226 , w6164 );
and ( w7228 , g47 , w6160 );
and ( w7229 , w7228 , g33 );
not ( w7230 , w7229 );
and ( w7231 , w7230 , w6136 );
and ( w7232 , w7227 , w7231 );
nor ( w7233 , w7232 , w7175 );
and ( w7234 , w7233 , w7263 );
not ( w7235 , w7234 );
and ( w7236 , w7235 , w6135 );
and ( w7237 , w7236 , w6134 );
and ( w7238 , w7237 , w6136 );
nor ( w7239 , w7238 , w6183 );
not ( w7240 , w7239 );
and ( w7241 , w7240 , w6136 );
nor ( w7242 , w7241 , w6785 );
not ( w7243 , w7242 );
and ( w7244 , w7243 , w6134 );
and ( w7245 , w7244 , w6791 );
and ( w7246 , w7245 , w6136 );
nor ( w7247 , w6797 , w7246 );
not ( w7248 , w7247 );
and ( w7249 , w7248 , w6135 );
and ( w7250 , w7249 , w6969 );
and ( w7251 , w7250 , w6135 );
and ( w7252 , w7251 , w6134 );
and ( w7253 , w7252 , w6136 );
and ( w7254 , w7253 , w6135 );
and ( w7255 , w7254 , w6791 );
and ( w7256 , w7255 , w6135 );
and ( w7257 , w7256 , w6134 );
nor ( w7258 , w6630 , w7257 );
not ( w7259 , w7258 );
and ( w7260 , w7259 , w6164 );
and ( w7261 , w7260 , w7231 );
nor ( w7262 , w7261 , w7175 );
not ( w7263 , w6878 );
and ( w7264 , w7262 , w7263 );
not ( w7265 , w7264 );
and ( w7266 , w7265 , w6135 );
and ( w7267 , w7266 , w6134 );
and ( w7268 , w7267 , w6136 );
nor ( w7269 , w7268 , w6183 );
not ( w7270 , w7269 );
and ( w7271 , w7270 , w6136 );
nor ( w7272 , w7271 , w6785 );
not ( w7273 , w7272 );
and ( w7274 , w7273 , w6791 );
and ( w7275 , w7274 , w6136 );
nor ( w7276 , w6605 , w7275 );
not ( w7277 , w7276 );
and ( w7278 , w7277 , w6136 );
and ( w7279 , w7278 , w6629 );
nor ( w7280 , w7279 , w7257 );
not ( w7281 , w7280 );
and ( w7282 , w7281 , w6136 );
and ( w7283 , w7282 , w6791 );
and ( w7284 , w7283 , w6135 );
and ( w7285 , w7284 , w6134 );
and ( w7286 , g39 , w7285 );
not ( w7287 , w7286 );
and ( w7288 , w7287 , w6160 );
and ( w7289 , g13 , w7285 );
not ( w7290 , w7289 );
and ( w7291 , w7288 , w7290 );
and ( w7292 , w7291 , w7354 );
not ( w7293 , w6193 );
and ( w7294 , w7293 , w7292 );
and ( w7295 , w7292 , w7356 );
and ( w7296 , w7285 , w7340 );
and ( w7297 , w7296 , w6169 );
and ( w7298 , w7297 , w7340 );
and ( w7299 , w7298 , w6134 );
and ( w7300 , w6606 , w7340 );
and ( w7301 , w7300 , w6136 );
and ( w7302 , w7301 , w6134 );
and ( w7303 , w7302 , w7285 );
and ( w7304 , w7299 , w7303 );
and ( w7305 , w7304 , w7297 );
and ( w7306 , w7305 , w7296 );
not ( w7307 , w7295 );
and ( w7308 , w7307 , w7306 );
and ( w7309 , w7308 , w7340 );
and ( w7310 , w7309 , w6134 );
and ( w7311 , w7310 , w6763 );
and ( w7312 , w7311 , w6969 );
and ( w7313 , w7285 , w6136 );
and ( w7314 , w7313 , w6169 );
and ( w7315 , w7314 , w6174 );
nor ( w7316 , w7315 , w6183 );
and ( w7317 , w7316 , w7292 );
not ( w7318 , w7317 );
and ( w7319 , w7318 , w6136 );
and ( w7320 , w7319 , w7340 );
and ( w7321 , w7320 , w6134 );
and ( w7322 , w7321 , w6135 );
and ( w7323 , w7322 , w6134 );
and ( w7324 , w7323 , w6177 );
and ( w7325 , w7324 , w6135 );
and ( w7326 , w7325 , w6878 );
nor ( w7327 , w7312 , w7326 );
and ( w7328 , w7294 , w7327 );
and ( w7329 , w7328 , w7348 );
and ( w7330 , w7327 , w7292 );
and ( w7331 , w7329 , w7330 );
and ( w7332 , w7331 , w7291 );
and ( w7333 , w7332 , w7327 );
not ( w7334 , w7333 );
and ( w7335 , w7334 , w7303 );
nor ( w7336 , w6763 , w7326 );
nor ( w7337 , w6133 , w7336 );
and ( w7338 , w7337 , w6134 );
and ( w7339 , w7335 , w7338 );
not ( w7340 , w6133 );
and ( w7341 , w7340 , w7339 );
and ( w7342 , w7341 , w6134 );
and ( w7343 , w6177 , w7342 );
and ( w7344 , w7350 , w7327 );
and ( w7345 , w7344 , w7292 );
and ( w7346 , w7345 , w7330 );
and ( w7347 , w7346 , w7327 );
not ( w7348 , w7326 );
and ( w7349 , w7344 , w7348 );
not ( w7350 , w7343 );
and ( w7351 , w7349 , w7350 );
and ( w7352 , w7347 , w7351 );
and ( w7353 , w7352 , w7291 );
not ( w7354 , w6183 );
and ( w7355 , w7353 , w7354 );
not ( w7356 , w6174 );
and ( w7357 , w7356 , w7355 );
not ( w7358 , w7357 );
and ( w7359 , w6169 , w7358 );
and ( w7360 , w6168 , w7359 );
and ( w7361 , w7360 , w7313 );
and ( w7362 , w6136 , w7339 );
and ( w7363 , w7361 , w7362 );
and ( w7364 , w7362 , w7313 );
not ( w7365 , w6629 );
and ( w7366 , w7365 , w7327 );
and ( w7367 , w7395 , w6134 );
and ( w7368 , w7367 , w6136 );
and ( w7369 , w7368 , w7395 );
and ( w7370 , w7364 , w7369 );
and ( w7371 , w7362 , w7369 );
and ( w7372 , w7370 , w7371 );
and ( w7373 , w7363 , w7372 );
and ( w7374 , w7373 , w7313 );
and ( w7375 , w7374 , w7369 );
nor ( w7376 , w6164 , w7375 );
not ( w7377 , w7376 );
and ( w7378 , w6136 , w7377 );
and ( w7379 , w7378 , w7313 );
and ( w7380 , w7379 , w7339 );
nor ( w7381 , w6133 , w7357 );
and ( w7382 , w7381 , w6134 );
and ( w7383 , w7380 , w7382 );
and ( w7384 , w7383 , w7359 );
and ( w7385 , w7384 , w7285 );
and ( w7386 , w7385 , w7313 );
and ( w7387 , w7386 , w7338 );
and ( w7388 , w6929 , w7382 );
and ( w7389 , w7388 , w7313 );
and ( w7390 , w7389 , w7369 );
and ( w7391 , w7390 , w7339 );
and ( w7392 , w7391 , w7372 );
and ( w7393 , w7392 , w7338 );
and ( w7394 , w7393 , w7369 );
not ( w7395 , w7366 );
and ( w7396 , w7394 , w7395 );
and ( w7397 , w7396 , w7359 );
nor ( w7398 , w7231 , w7397 );
not ( w7399 , w7398 );
and ( t_1 , w7387 , w7399 );
and ( w7400 , w12921 , w485 );
and ( w7401 , w7400 , w105 );
not ( w7402 , w73 );
and ( w7403 , w7402 , g5 );
not ( w7404 , w7403 );
and ( w7405 , w7404 , g5 );
not ( w7406 , w7405 );
and ( w7407 , w11 , w7406 );
not ( w7408 , w7407 );
and ( w7409 , w7408 , g5 );
and ( w7410 , w11092 , w52 );
nor ( w7411 , w7409 , w7410 );
and ( w7412 , g6 , w12934 );
and ( w7413 , w7412 , w11092 );
nor ( w7414 , w222 , w7413 );
not ( w7415 , w224 );
and ( w7416 , w7414 , w7415 );
nor ( w7417 , w1 , w7416 );
nor ( w7418 , w7417 , w7413 );
not ( w7419 , w212 );
and ( w7420 , w7419 , w7418 );
nor ( w7421 , w11 , w8 );
nor ( w7422 , w7421 , w2551 );
nor ( w7423 , w7422 , g5 );
nor ( w7424 , w7423 , w7409 );
nor ( w7425 , w7420 , w7424 );
not ( w7426 , w206 );
and ( w7427 , w7426 , g7 );
nor ( w7428 , w7427 , w7405 );
not ( w7429 , w7425 );
and ( w7430 , w7429 , w7428 );
and ( w7431 , w7411 , w7430 );
and ( w7432 , w7431 , w7418 );
nor ( w7433 , w7432 , w7424 );
not ( w7434 , w7433 );
and ( w7435 , w7434 , w7428 );
not ( w7436 , w4 );
and ( w7437 , w7436 , g5 );
not ( w7438 , w2728 );
and ( w7439 , w7438 , g7 );
nor ( w7440 , w7439 , g6 );
nor ( w7441 , w7440 , g6 );
nor ( w7442 , w69 , w2623 );
not ( w7443 , w7441 );
and ( w7444 , w7443 , w7442 );
and ( w7445 , w7444 , w7457 );
not ( w7446 , w7437 );
and ( w7447 , w7446 , w7445 );
and ( w7448 , w7418 , w7447 );
and ( w7449 , w7435 , w7448 );
nor ( w7450 , w7449 , w43 );
and ( w7451 , w13206 , w7428 );
nor ( w7452 , g31 , w7451 );
nor ( w7453 , w7450 , w7452 );
nor ( w7454 , w8 , g7 );
and ( w7455 , w7454 , w11092 );
nor ( w7456 , w7439 , w7455 );
not ( w7457 , w2623 );
and ( w7458 , w7456 , w7457 );
and ( w7459 , w7458 , w7428 );
and ( w7460 , w7453 , w7459 );
and ( w7461 , w7460 , w12919 );
nor ( w7462 , w7461 , w7449 );
nor ( w7463 , w7462 , w485 );
nor ( w7464 , w7463 , w48 );
not ( w7465 , w7464 );
and ( w7466 , w7465 , w7428 );
nor ( w7467 , w7466 , w20 );
not ( w7468 , w21 );
and ( w7469 , w7468 , g15 );
and ( w7470 , w7469 , g14 );
not ( w7471 , w7470 );
and ( w7472 , w7471 , g14 );
and ( w7473 , w7472 , g15 );
and ( w7474 , w7473 , g17 );
nor ( w7475 , w7474 , g16 );
nor ( w7476 , w56 , w21 );
and ( w7477 , w7476 , g16 );
and ( w7478 , w7477 , w7445 );
and ( w7479 , w7478 , w7458 );
nor ( w7480 , w7475 , w7479 );
nor ( w7481 , w7480 , w272 );
and ( w7482 , w7481 , w7445 );
and ( w7483 , w7482 , w7458 );
nor ( w7484 , w274 , w7483 );
not ( w7485 , w31 );
and ( w7486 , w7484 , w7485 );
and ( w7487 , w7499 , w7459 );
nor ( w7488 , w7487 , w37 );
not ( w7489 , w7488 );
and ( w7490 , w7489 , w7459 );
nor ( w7491 , w7490 , w41 );
nor ( w7492 , w7491 , w39 );
and ( w7493 , w7492 , w7459 );
and ( w7494 , w9049 , g16 );
nor ( w7495 , w56 , w7494 );
and ( w7496 , g16 , w7495 );
nor ( w7497 , w33 , w7496 );
and ( w7498 , w7497 , w11140 );
not ( w7499 , w7486 );
and ( w7500 , w7499 , w7498 );
and ( w7501 , w7500 , w8363 );
nor ( w7502 , w7501 , w37 );
nor ( w7503 , w7502 , w39 );
and ( w7504 , w7503 , w7445 );
nor ( w7505 , w41 , w7504 );
not ( w7506 , w7505 );
and ( w7507 , w7506 , w7445 );
and ( w7508 , w7493 , w7507 );
and ( w7509 , w7508 , w7459 );
and ( w7510 , w7509 , w12117 );
and ( w7511 , w7510 , w7458 );
and ( w7512 , w7511 , w7428 );
and ( w7513 , w7512 , w7448 );
nor ( w7514 , w7513 , w43 );
and ( w7515 , w12117 , w41 );
nor ( w7516 , w7515 , w43 );
and ( w7517 , w7516 , w12142 );
not ( w7518 , w7517 );
and ( w7519 , w7518 , w7428 );
nor ( w7520 , w7519 , w7435 );
not ( w7521 , w7520 );
and ( w7522 , w7521 , w7428 );
not ( w7523 , w7522 );
and ( w7524 , w7514 , w7523 );
and ( w7525 , w485 , w18 );
not ( w7526 , w7525 );
and ( w7527 , w7526 , w7448 );
not ( w7528 , w7524 );
and ( w7529 , w7528 , w7527 );
not ( w7530 , w7529 );
and ( w7531 , w7530 , w485 );
nor ( w7532 , w7514 , w7452 );
and ( w7533 , w7532 , w7459 );
and ( w7534 , w7533 , w12919 );
nor ( w7535 , w7534 , w48 );
not ( w7536 , w7535 );
and ( w7537 , w7536 , w7458 );
and ( w7538 , w7537 , w7428 );
and ( w7539 , w7538 , w7448 );
nor ( w7540 , w7539 , w485 );
not ( w7541 , w7540 );
and ( w7542 , w7541 , w7448 );
not ( w7543 , w7531 );
and ( w7544 , w7543 , w7542 );
nor ( w7545 , w7544 , w48 );
and ( w7546 , w7545 , w12921 );
and ( w7547 , w7546 , w11166 );
and ( w7548 , w255 , w7428 );
and ( w7549 , w7548 , w7448 );
not ( w7550 , w7549 );
and ( w7551 , w7547 , w7550 );
and ( w7552 , w7551 , w8876 );
not ( w7553 , w7552 );
and ( w7554 , w7553 , w7428 );
and ( w7555 , w7554 , w7448 );
and ( w7556 , w7467 , w8829 );
and ( w7557 , w7556 , w8848 );
nor ( w7558 , w377 , g28 );
and ( w7559 , w7558 , w13333 );
nor ( w7560 , w7559 , g31 );
and ( w7561 , w7560 , w7458 );
and ( w7562 , w7561 , w7428 );
nor ( w7563 , w7562 , g31 );
not ( w7564 , w4430 );
and ( w7565 , w7564 , g31 );
not ( w7566 , w7565 );
and ( w7567 , w7566 , w310 );
nor ( w7568 , w7567 , w7435 );
and ( w7569 , w7568 , w8272 );
not ( w7570 , w7569 );
and ( w7571 , w7570 , w7458 );
and ( w7572 , w7571 , w7428 );
and ( w7573 , w7572 , g30 );
not ( w7574 , w7573 );
and ( w7575 , w7574 , g30 );
not ( w7576 , w7575 );
and ( w7577 , w7576 , g31 );
not ( w7578 , w7577 );
and ( w7579 , w7578 , g31 );
not ( w7580 , w7579 );
and ( w7581 , w7580 , w7458 );
nor ( w7582 , w7581 , w7435 );
not ( w7583 , w7582 );
and ( w7584 , w7583 , w7428 );
and ( w7585 , w7584 , w7448 );
not ( w7586 , w7563 );
and ( w7587 , w7586 , w7585 );
and ( w7588 , w7587 , w7459 );
nor ( w7589 , w7561 , g31 );
and ( w7590 , w7618 , w7459 );
and ( w7591 , w7590 , w7458 );
and ( w7592 , w7591 , w7428 );
and ( w7593 , w7588 , w7592 );
and ( w7594 , w7593 , w7458 );
and ( w7595 , w7594 , w7428 );
and ( w7596 , w7595 , w7418 );
and ( w7597 , w7596 , w7448 );
nor ( w7598 , w7449 , w7513 );
and ( w7599 , w7598 , w12144 );
and ( w7600 , w7599 , w12919 );
and ( w7601 , w12919 , w7459 );
and ( w7602 , w7601 , w7458 );
nor ( w7603 , w7602 , w7435 );
not ( w7604 , w7603 );
and ( w7605 , w7604 , w7428 );
and ( w7606 , w7605 , w7448 );
not ( w7607 , w7600 );
and ( w7608 , w7607 , w7606 );
and ( w7609 , w7428 , w7585 );
and ( w7610 , w7609 , w7459 );
and ( w7611 , w7610 , w7592 );
and ( w7612 , w7611 , w7458 );
and ( w7613 , w7612 , w7428 );
and ( w7614 , w7613 , w7418 );
and ( w7615 , w7614 , w7448 );
and ( w7616 , w7618 , w7615 );
and ( w7617 , w7616 , w43 );
not ( w7618 , w7589 );
and ( w7619 , w7618 , w7428 );
and ( w7620 , w7619 , w7585 );
and ( w7621 , w7620 , w7459 );
and ( w7622 , w7621 , w7592 );
nor ( w7623 , w274 , w31 );
and ( w7624 , w7504 , w11140 );
and ( w7625 , w7624 , w7418 );
and ( w7626 , w7625 , w7458 );
and ( w7627 , w7817 , w7626 );
and ( w7628 , w7627 , w8363 );
and ( w7629 , w7627 , w7418 );
nor ( w7630 , w7629 , w7424 );
not ( w7631 , w7630 );
and ( w7632 , w7631 , w7458 );
and ( w7633 , w7632 , w7428 );
and ( w7634 , w7628 , w7633 );
not ( w7635 , w429 );
and ( w7636 , w7635 , w7418 );
not ( w7637 , w7636 );
and ( w7638 , w21 , w7637 );
nor ( w7639 , w7638 , w56 );
and ( w7640 , w7639 , w7418 );
not ( w7641 , w7640 );
and ( w7642 , w21 , w7641 );
nor ( w7643 , w7642 , w56 );
and ( w7644 , w7643 , w8363 );
and ( w7645 , w7644 , w11347 );
and ( w7646 , w31 , w7633 );
nor ( w7647 , w7646 , w7483 );
and ( w7648 , w7647 , g19 );
not ( w7649 , w7648 );
and ( w7650 , w7649 , w7418 );
nor ( w7651 , w7650 , w7424 );
not ( w7652 , w7651 );
and ( w7653 , w7652 , w7458 );
and ( w7654 , w7653 , w7428 );
and ( w7655 , w7645 , w7654 );
and ( w7656 , w7655 , w11140 );
nor ( w7657 , w7656 , w7435 );
not ( w7658 , w7657 );
and ( w7659 , w7658 , w7418 );
nor ( w7660 , w7659 , w7424 );
not ( w7661 , w7660 );
and ( w7662 , w7661 , w7458 );
and ( w7663 , w7662 , w7428 );
nor ( w7664 , w7634 , w7663 );
and ( w7665 , w7664 , w12424 );
and ( w7666 , w7665 , w7803 );
not ( w7667 , w7666 );
and ( w7668 , w7667 , w7458 );
and ( w7669 , w7668 , w7428 );
and ( w7670 , w7669 , w7418 );
and ( w7671 , w7670 , w7448 );
and ( w7672 , w7622 , w7671 );
not ( w7673 , w7496 );
and ( w7674 , w7672 , w7673 );
nor ( w7675 , w7674 , w48 );
not ( w7676 , w7675 );
and ( w7677 , w7676 , w7459 );
and ( w7678 , w7677 , w7458 );
and ( w7679 , w7678 , w7428 );
and ( w7680 , w7679 , w7418 );
and ( w7681 , w7680 , w7448 );
and ( w7682 , w12144 , w7681 );
nor ( w7683 , w7682 , w7435 );
not ( w7684 , w7683 );
and ( w7685 , w7684 , w7448 );
nor ( w7686 , w7617 , w7685 );
not ( w7687 , w7686 );
and ( w7688 , w7687 , w7458 );
and ( w7689 , w7688 , w7428 );
and ( w7690 , w7689 , w7418 );
and ( w7691 , w7690 , w7448 );
not ( w7692 , w7691 );
and ( w7693 , w7450 , w7692 );
and ( w7694 , w7693 , w12717 );
nor ( w7695 , w7694 , w18 );
and ( w7696 , w7695 , w7615 );
and ( w7697 , w7696 , w7585 );
nor ( w7698 , w7697 , w18 );
and ( w7699 , w12919 , w7496 );
not ( w7700 , w7699 );
and ( w7701 , w7700 , w7458 );
and ( w7702 , w7701 , w7428 );
and ( w7703 , w7702 , w7448 );
not ( w7704 , w7698 );
and ( w7705 , w7704 , w7703 );
nor ( w7706 , w7705 , w20 );
and ( w7707 , w7706 , w12142 );
not ( w7708 , w7707 );
and ( w7709 , w7708 , w7428 );
and ( w7710 , w7709 , w11852 );
and ( w7711 , w7710 , w7459 );
and ( w7712 , w3577 , w7448 );
and ( w7713 , w7711 , w7712 );
nor ( w7714 , w7515 , w7435 );
not ( w7715 , w7714 );
and ( w7716 , w7715 , w7428 );
nor ( w7717 , w7716 , w7513 );
nor ( w7718 , w43 , w48 );
not ( w7719 , w7718 );
and ( w7720 , w7719 , w7428 );
nor ( w7721 , w7720 , w7435 );
not ( w7722 , w7721 );
and ( w7723 , w7722 , w7428 );
and ( w7724 , w7717 , w7773 );
and ( w7725 , w7724 , w12144 );
nor ( w7726 , w7725 , w18 );
and ( w7727 , w7726 , w7527 );
nor ( w7728 , w7727 , w48 );
and ( w7729 , w7728 , w12921 );
and ( w7730 , w7729 , w485 );
not ( w7731 , w7514 );
and ( w7732 , w7731 , w7459 );
and ( w7733 , w7732 , w12919 );
nor ( w7734 , w7733 , w48 );
and ( w7735 , w7734 , w12921 );
and ( w7736 , w7735 , w8640 );
not ( w7737 , w7736 );
and ( w7738 , w7737 , w7458 );
and ( w7739 , w7738 , w7428 );
and ( w7740 , w7739 , w7448 );
not ( w7741 , w7730 );
and ( w7742 , w7741 , w7740 );
nor ( w7743 , w7742 , w105 );
and ( w7744 , g32 , w13211 );
and ( w7745 , g32 , w8002 );
and ( w7746 , w7745 , w7448 );
not ( w7747 , w7746 );
and ( w7748 , w7743 , w7747 );
and ( w7749 , w7748 , w255 );
and ( w7750 , w7749 , w8876 );
not ( w7751 , w7750 );
and ( w7752 , w7751 , w7428 );
and ( w7753 , w7752 , w7448 );
and ( w7754 , w8845 , w7753 );
nor ( w7755 , w7754 , w7746 );
and ( w7756 , w7755 , w8848 );
not ( w7757 , w7756 );
and ( w7758 , w7757 , w7712 );
and ( w7759 , w7758 , w8848 );
and ( w7760 , w485 , w8848 );
nor ( w7761 , w5252 , w7760 );
and ( w7762 , w7759 , w8036 );
not ( w7763 , w7762 );
and ( w7764 , w7763 , w255 );
and ( w7765 , w8845 , w7555 );
nor ( w7766 , w7765 , w7746 );
not ( w7767 , w7766 );
and ( w7768 , w7767 , w7712 );
and ( w7769 , w7768 , w8036 );
and ( w7770 , w8848 , w7769 );
nor ( w7771 , w7770 , w7549 );
and ( w7772 , w7717 , w12144 );
not ( w7773 , w7723 );
and ( w7774 , w7772 , w7773 );
nor ( w7775 , w7774 , w18 );
and ( w7776 , w7775 , w7527 );
nor ( w7777 , w7776 , w48 );
and ( w7778 , w7777 , w12921 );
and ( w7779 , w7778 , w485 );
and ( w7780 , w7514 , w12919 );
nor ( w7781 , w7601 , w7449 );
nor ( w7782 , w7716 , w7723 );
and ( w7783 , w7782 , w8305 );
and ( w7784 , w7783 , w12144 );
not ( w7785 , w7784 );
and ( w7786 , w7785 , w7527 );
nor ( w7787 , w7786 , w48 );
and ( w7788 , w7787 , w12921 );
and ( w7789 , w7788 , w485 );
and ( w7790 , w11226 , g33 );
nor ( w7791 , w7790 , w7744 );
and ( w7792 , w7791 , w7458 );
and ( w7793 , w7792 , w7428 );
and ( w7794 , w7459 , w7793 );
not ( w7795 , w7483 );
and ( w7796 , w7623 , w7795 );
not ( w7797 , w7796 );
and ( w7798 , w7797 , w7498 );
and ( w7799 , w7798 , w8363 );
nor ( w7800 , w7799 , w37 );
nor ( w7801 , w7800 , w39 );
nor ( w7802 , w7801 , w43 );
not ( w7803 , w41 );
and ( w7804 , w7802 , w7803 );
nor ( w7805 , w7804 , w45 );
nor ( w7806 , w7805 , w48 );
nor ( w7807 , w7806 , w105 );
and ( w7808 , w7807 , w12919 );
and ( w7809 , w7808 , w7445 );
and ( w7810 , w7809 , w7458 );
and ( w7811 , w7794 , w7810 );
and ( w7812 , w8640 , w105 );
nor ( w7813 , w7812 , w19 );
nor ( w7814 , w7811 , w7813 );
and ( w7815 , w7814 , w12498 );
nor ( w7816 , w7720 , w7810 );
not ( w7817 , w7623 );
and ( w7818 , w7817 , w7633 );
and ( w7819 , w7818 , w7626 );
nor ( w7820 , w7819 , w43 );
and ( w7821 , w7820 , w12142 );
and ( w7822 , w7459 , w7418 );
nor ( w7823 , w7822 , w7424 );
not ( w7824 , w7823 );
and ( w7825 , w7824 , w7428 );
not ( w7826 , w7821 );
and ( w7827 , w7826 , w7825 );
nor ( w7828 , w7827 , w7435 );
not ( w7829 , w7828 );
and ( w7830 , w7829 , w7418 );
nor ( w7831 , w7830 , w7424 );
not ( w7832 , w7831 );
and ( w7833 , w7832 , w7458 );
and ( w7834 , w7833 , w7428 );
and ( w7835 , w7880 , w7834 );
and ( w7836 , w35 , w8876 );
and ( w7837 , w7835 , w7907 );
nor ( w7838 , w7663 , w7435 );
and ( w7839 , w7838 , w12144 );
and ( w7840 , w7839 , w12142 );
not ( w7841 , w7840 );
and ( w7842 , w7841 , w7825 );
and ( w7843 , w7459 , w7418 );
nor ( w7844 , w7843 , w7424 );
not ( w7845 , w7844 );
and ( w7846 , w7845 , w7458 );
and ( w7847 , w7846 , w7428 );
and ( w7848 , w7842 , w7847 );
and ( w7849 , w7848 , w7459 );
and ( w7850 , w7849 , w12919 );
nor ( w7851 , w7850 , w7435 );
not ( w7852 , w7851 );
and ( w7853 , w7852 , w7418 );
nor ( w7854 , w7853 , w7424 );
not ( w7855 , w7854 );
and ( w7856 , w7855 , w7458 );
and ( w7857 , w7856 , w7428 );
and ( w7858 , w7880 , w7857 );
and ( w7859 , w7858 , w12919 );
nor ( w7860 , w7859 , w7435 );
and ( w7861 , w7860 , w8272 );
not ( w7862 , w7861 );
and ( w7863 , w7862 , w7458 );
and ( w7864 , w7863 , w11166 );
and ( w7865 , w7864 , w7428 );
nor ( w7866 , w7837 , w7865 );
nor ( w7867 , w37 , w41 );
nor ( w7868 , w7867 , w39 );
nor ( w7869 , w7868 , w43 );
and ( w7870 , w7869 , w12142 );
not ( w7871 , w7870 );
and ( w7872 , w7871 , w7825 );
nor ( w7873 , w7872 , w7435 );
not ( w7874 , w7873 );
and ( w7875 , w7874 , w7418 );
nor ( w7876 , w7875 , w7424 );
not ( w7877 , w7876 );
and ( w7878 , w7877 , w7458 );
and ( w7879 , w7878 , w7428 );
not ( w7880 , w7816 );
and ( w7881 , w7880 , w7879 );
nor ( w7882 , w7881 , w20 );
nor ( w7883 , w7882 , w18 );
nor ( w7884 , w7883 , w7435 );
not ( w7885 , w7884 );
and ( w7886 , w7885 , w7418 );
nor ( w7887 , w7886 , w7424 );
not ( w7888 , w7887 );
and ( w7889 , w7888 , w7458 );
and ( w7890 , w7889 , w11166 );
and ( w7891 , w7890 , w7428 );
not ( w7892 , w7891 );
and ( w7893 , w7866 , w7892 );
and ( w7894 , w7893 , w12921 );
not ( w7895 , w7894 );
and ( w7896 , w7895 , w7847 );
and ( w7897 , w7896 , w8002 );
and ( w7898 , w7897 , w12037 );
and ( w7899 , w7898 , w13211 );
and ( w7900 , w48 , w7428 );
nor ( w7901 , w7900 , w43 );
nor ( w7902 , w7901 , w18 );
nor ( w7903 , w7902 , w7810 );
not ( w7904 , w7818 );
and ( w7905 , w7904 , w7838 );
nor ( w7906 , w7905 , w33 );
not ( w7907 , w7836 );
and ( w7908 , w7906 , w7907 );
nor ( w7909 , w7908 , w37 );
nor ( w7910 , w7909 , w39 );
nor ( w7911 , w7910 , w41 );
and ( w7912 , w7911 , w12142 );
and ( w7913 , w7912 , w12717 );
and ( w7914 , w7913 , w12144 );
and ( w7915 , w7914 , w8876 );
not ( w7916 , w7915 );
and ( w7917 , w7916 , w7418 );
nor ( w7918 , w7917 , w7424 );
not ( w7919 , w7918 );
and ( w7920 , w7919 , w7458 );
and ( w7921 , w7920 , w7428 );
and ( w7922 , w7458 , w7921 );
nor ( w7923 , w18 , w7922 );
not ( w7924 , w7479 );
and ( w7925 , g16 , w7924 );
nor ( w7926 , w7925 , g17 );
and ( w7927 , w21 , w9049 );
nor ( w7928 , w7927 , w7424 );
not ( w7929 , w7928 );
and ( w7930 , w7929 , w7458 );
and ( w7931 , w7930 , w7428 );
nor ( w7932 , w7926 , w7931 );
and ( w7933 , w7932 , w8272 );
not ( w7934 , w7933 );
and ( w7935 , w7934 , w7428 );
nor ( w7936 , g17 , w7935 );
not ( w7937 , w7936 );
and ( w7938 , w7937 , w7459 );
and ( w7939 , w7938 , w7458 );
and ( w7940 , w7939 , w7428 );
not ( w7941 , w7923 );
and ( w7942 , w7941 , w7940 );
and ( w7943 , w7942 , w7418 );
nor ( w7944 , w7943 , w7424 );
not ( w7945 , w7944 );
and ( w7946 , w7945 , w7458 );
and ( w7947 , w7946 , w7428 );
not ( w7948 , w7903 );
and ( w7949 , w7948 , w7947 );
nor ( w7950 , w7949 , w20 );
not ( w7951 , w7950 );
and ( w7952 , w7951 , w7847 );
not ( w7953 , w7952 );
and ( w7954 , w7953 , w312 );
and ( w7955 , w7954 , w8876 );
not ( w7956 , w7955 );
and ( w7957 , w7956 , w7418 );
nor ( w7958 , w7957 , w7424 );
not ( w7959 , w7958 );
and ( w7960 , w7959 , w7458 );
and ( w7961 , w7960 , w11166 );
and ( w7962 , w7961 , w7428 );
and ( w7963 , g32 , w7962 );
and ( w7964 , w7963 , w7459 );
and ( w7965 , w7964 , w12532 );
and ( w7966 , w7965 , g33 );
nor ( w7967 , w7966 , w7435 );
not ( w7968 , w7967 );
and ( w7969 , w7968 , w7458 );
and ( w7970 , w7969 , w7428 );
nor ( w7971 , w7899 , w7970 );
nor ( w7972 , w7971 , w18 );
and ( w7973 , w7810 , w7572 );
nor ( w7974 , w7973 , w7435 );
and ( w7975 , w7974 , w8272 );
not ( w7976 , w7975 );
and ( w7977 , w7976 , w7428 );
nor ( w7978 , w7972 , w7977 );
and ( w7979 , w7978 , w8876 );
not ( w7980 , w7979 );
and ( w7981 , w7980 , w7418 );
nor ( w7982 , w7981 , w7424 );
not ( w7983 , w7982 );
and ( w7984 , w7983 , w7458 );
and ( w7985 , w7984 , w11166 );
and ( w7986 , w7985 , w7428 );
and ( w7987 , w7794 , w7986 );
nor ( w7988 , w7987 , g28 );
and ( w7989 , w7988 , w13333 );
not ( w7990 , w7989 );
and ( w7991 , w7990 , w7459 );
and ( w7992 , w7459 , w7810 );
nor ( w7993 , w7992 , w7813 );
and ( w7994 , w7993 , w12498 );
and ( w7995 , w7994 , w19 );
and ( w7996 , w7995 , w8272 );
not ( w7997 , w7996 );
and ( w7998 , w7997 , w7458 );
and ( w7999 , w7998 , w11166 );
and ( w8000 , w7999 , w7428 );
and ( w8001 , w7991 , w8000 );
not ( w8002 , w7744 );
and ( w8003 , w8002 , w7458 );
and ( w8004 , w8003 , w7428 );
not ( w8005 , w7790 );
and ( w8006 , w8005 , w8004 );
and ( w8007 , w8006 , w7459 );
and ( w8008 , w8001 , w8007 );
nor ( w8009 , w8008 , w7435 );
not ( w8010 , w8009 );
and ( w8011 , w8010 , w19 );
and ( w8012 , w8011 , w7418 );
not ( w8013 , w8012 );
and ( w8014 , w8013 , w19 );
and ( w8015 , w8014 , w8272 );
not ( w8016 , w8015 );
and ( w8017 , w8016 , w7458 );
and ( w8018 , w8017 , w11166 );
and ( w8019 , w8018 , w7428 );
not ( w8020 , w7815 );
and ( w8021 , w8020 , w8019 );
and ( w8022 , w8021 , w8007 );
not ( w8023 , w8022 );
and ( w8024 , w8023 , w19 );
and ( w8025 , w8024 , w8272 );
not ( w8026 , w8025 );
and ( w8027 , w8026 , w7458 );
and ( w8028 , w8027 , w11166 );
and ( w8029 , w8028 , w7428 );
and ( w8030 , w19 , w8029 );
and ( w8031 , w8030 , w7458 );
and ( w8032 , w8031 , w7428 );
and ( w8033 , w8032 , w7418 );
and ( w8034 , w8033 , w7448 );
nor ( w8035 , w8034 , w19 );
not ( w8036 , w7761 );
and ( w8037 , w8036 , w7448 );
nor ( w8038 , w7813 , w7435 );
and ( w8039 , w8636 , w8038 );
not ( w8040 , w8039 );
and ( w8041 , w8040 , w7448 );
nor ( w8042 , w7449 , w8041 );
not ( w8043 , w7813 );
and ( w8044 , w8042 , w8043 );
nor ( w8045 , w20 , g10 );
and ( w8046 , w8045 , w105 );
not ( w8047 , w8046 );
and ( w8048 , w8047 , g11 );
and ( w8049 , w12921 , w105 );
nor ( w8050 , w8049 , w19 );
nor ( w8051 , w8050 , w7760 );
not ( w8052 , w8048 );
and ( w8053 , w8052 , w8051 );
and ( w8054 , w8053 , w8798 );
not ( w8055 , w8054 );
and ( w8056 , w8055 , w7445 );
and ( w8057 , w8056 , w7458 );
and ( w8058 , w8848 , w8057 );
and ( w8059 , w8058 , w7428 );
and ( w8060 , w8059 , w7448 );
and ( w8061 , w8044 , w8634 );
not ( w8062 , w8029 );
and ( w8063 , w8061 , w8062 );
and ( w8064 , w8063 , w8594 );
and ( w8065 , w8064 , w8798 );
and ( w8066 , w8065 , w8876 );
not ( w8067 , w8066 );
and ( w8068 , w8067 , w7448 );
not ( w8069 , w8035 );
and ( w8070 , w8069 , w8068 );
and ( w8071 , w8070 , w7458 );
and ( w8072 , w8071 , w7428 );
and ( w8073 , w8072 , w7418 );
and ( w8074 , w8073 , w7448 );
nor ( w8075 , w7733 , w8074 );
and ( w8076 , w8075 , w12142 );
and ( w8077 , w8076 , w12921 );
and ( w8078 , w8077 , w8640 );
and ( w8079 , w8078 , w12498 );
not ( w8080 , w8079 );
and ( w8081 , w8080 , w7459 );
not ( w8082 , w7484 );
and ( w8083 , w8082 , w7459 );
nor ( w8084 , w8083 , w31 );
not ( w8085 , w8084 );
and ( w8086 , w8085 , w7459 );
nor ( w8087 , w8086 , w37 );
not ( w8088 , w8087 );
and ( w8089 , w8088 , w7459 );
nor ( w8090 , w8089 , w41 );
nor ( w8091 , w8090 , w39 );
and ( w8092 , w8091 , w7459 );
and ( w8093 , w8092 , w7507 );
and ( w8094 , w8093 , w7459 );
and ( w8095 , w8094 , w12117 );
nor ( w8096 , w8095 , w7449 );
and ( w8097 , w8096 , w12919 );
not ( w8098 , w8097 );
and ( w8099 , w8098 , w7458 );
nor ( w8100 , w8099 , w7435 );
not ( w8101 , w8100 );
and ( w8102 , w8101 , w7428 );
and ( w8103 , w8102 , w7448 );
and ( w8104 , w12919 , w8103 );
nor ( w8105 , w8104 , w48 );
nor ( w8106 , g33 , w7744 );
nor ( w8107 , w8106 , w7746 );
not ( w8108 , w8107 );
and ( w8109 , w8108 , w7448 );
not ( w8110 , w8105 );
and ( w8111 , w8110 , w8109 );
nor ( w8112 , w8041 , w8060 );
not ( w8113 , w8112 );
and ( w8114 , w8113 , w105 );
and ( w8115 , w7601 , w8103 );
nor ( w8116 , w8115 , w48 );
not ( w8117 , w8116 );
and ( w8118 , w8117 , w7428 );
nor ( w8119 , w8118 , w20 );
not ( w8120 , w8119 );
and ( w8121 , w8120 , w7459 );
and ( w8122 , w8121 , w377 );
nor ( w8123 , w8089 , w41 );
not ( w8124 , w8123 );
and ( w8125 , w8124 , w7459 );
nor ( w8126 , w384 , w7435 );
not ( w8127 , w8126 );
and ( w8128 , w8125 , w8127 );
and ( w8129 , w8125 , w7507 );
and ( w8130 , w8129 , w7458 );
and ( w8131 , w8130 , w7428 );
and ( w8132 , w8131 , w7448 );
and ( w8133 , w8132 , w11852 );
nor ( w8134 , w8133 , w20 );
and ( w8135 , w8134 , w8640 );
not ( w8136 , w8135 );
and ( w8137 , w8136 , w7448 );
nor ( w8138 , w8128 , w8137 );
not ( w8139 , w8138 );
and ( w8140 , w8139 , w7459 );
and ( w8141 , w8140 , w11140 );
and ( w8142 , w8141 , w7507 );
and ( w8143 , w8142 , w7459 );
and ( w8144 , w8143 , w12117 );
and ( w8145 , w8144 , w7459 );
and ( w8146 , w8145 , w12919 );
nor ( w8147 , w8146 , w20 );
not ( w8148 , w8147 );
and ( w8149 , w8148 , w7458 );
nor ( w8150 , w8149 , w7435 );
not ( w8151 , w8150 );
and ( w8152 , w8151 , w7428 );
and ( w8153 , w8152 , w7448 );
nor ( w8154 , w48 , w8153 );
and ( w8155 , w8154 , w12919 );
not ( w8156 , w8155 );
and ( w8157 , w8156 , w7459 );
and ( w8158 , w8157 , w12919 );
nor ( w8159 , w8158 , w8034 );
nor ( w8160 , w20 , w8159 );
nor ( w8161 , w8160 , w19 );
not ( w8162 , w8161 );
and ( w8163 , w8162 , w8029 );
and ( w8164 , w8163 , w11166 );
and ( w8165 , w8640 , w8164 );
and ( w8166 , w8165 , w12080 );
and ( w8167 , w8166 , w7458 );
and ( w8168 , w8167 , w7428 );
and ( w8169 , w8168 , w7418 );
and ( w8170 , w8169 , w7448 );
nor ( w8171 , w8122 , w8170 );
and ( w8172 , w8171 , w8848 );
not ( w8173 , w8172 );
and ( w8174 , w8173 , w8029 );
and ( w8175 , w8174 , w11166 );
nor ( w8176 , w8175 , w485 );
and ( w8177 , w8176 , w8247 );
nor ( w8178 , w8177 , w485 );
and ( w8179 , w8178 , w12080 );
and ( w8180 , w8179 , w7458 );
nor ( w8181 , w8180 , w7435 );
not ( w8182 , w8181 );
and ( w8183 , w8182 , w7428 );
and ( w8184 , w8183 , w7418 );
and ( w8185 , w8184 , w7448 );
nor ( w8186 , w8114 , w8185 );
and ( w8187 , w8186 , w8640 );
and ( w8188 , w8187 , w8247 );
nor ( w8189 , w8188 , w485 );
nor ( w8190 , w8189 , w7435 );
not ( w8191 , w8190 );
and ( w8192 , w8191 , w7428 );
and ( w8193 , w8192 , w7448 );
and ( w8194 , w8111 , w8193 );
and ( w8195 , w8194 , w7459 );
and ( w8196 , w8195 , w377 );
nor ( w8197 , w8196 , w8074 );
and ( w8198 , w8197 , w12921 );
and ( w8199 , w8198 , w8640 );
and ( w8200 , w8199 , w8247 );
nor ( w8201 , w8200 , w485 );
and ( w8202 , w8201 , w11166 );
nor ( w8203 , w8202 , w19 );
not ( w8204 , w8203 );
and ( w8205 , w8204 , w8068 );
and ( w8206 , w8205 , w7458 );
nor ( w8207 , w8206 , w7435 );
not ( w8208 , w8207 );
and ( w8209 , w8208 , w7428 );
and ( w8210 , w8209 , w7418 );
and ( w8211 , w8210 , w7448 );
nor ( w8212 , w8211 , w7527 );
and ( w8213 , w8212 , w485 );
not ( w8214 , w7810 );
and ( w8215 , w8213 , w8214 );
not ( w8216 , w8215 );
and ( w8217 , w8216 , w485 );
nor ( w8218 , w8211 , w48 );
and ( w8219 , w8218 , w18 );
not ( w8220 , w8219 );
and ( w8221 , w8220 , w7459 );
nor ( w8222 , w8221 , w20 );
and ( w8223 , w7514 , w12142 );
and ( w8224 , w8223 , w12919 );
nor ( w8225 , w20 , w8074 );
and ( w8226 , w8225 , w8640 );
nor ( w8227 , w8226 , w105 );
and ( w8228 , w8227 , w8068 );
and ( w8229 , w8228 , w7448 );
not ( w8230 , w8229 );
and ( w8231 , w8224 , w8230 );
and ( w8232 , w8231 , w12498 );
not ( w8233 , w8232 );
and ( w8234 , w8233 , w7459 );
nor ( w8235 , w8234 , w485 );
and ( w8236 , w8235 , w12921 );
and ( w8237 , w7450 , w12142 );
nor ( w8238 , w8237 , w18 );
nor ( w8239 , w8238 , w48 );
not ( w8240 , w8239 );
and ( w8241 , w8240 , w7428 );
and ( w8242 , w8241 , w7459 );
and ( w8243 , w8242 , w377 );
nor ( w8244 , w8243 , w8034 );
nor ( w8245 , w20 , w8244 );
nor ( w8246 , w8245 , w485 );
not ( w8247 , w7449 );
and ( w8248 , w8246 , w8247 );
nor ( w8249 , w8248 , w485 );
nor ( w8250 , w8249 , w19 );
not ( w8251 , w8250 );
and ( w8252 , w8251 , w8029 );
and ( w8253 , w8252 , w11166 );
and ( w8254 , w8253 , w7458 );
nor ( w8255 , w8254 , w7435 );
not ( w8256 , w8255 );
and ( w8257 , w8256 , w7428 );
and ( w8258 , w8257 , w7418 );
and ( w8259 , w8258 , w7448 );
nor ( w8260 , w8259 , w8229 );
nor ( w8261 , w310 , g30 );
and ( w8262 , w8261 , g31 );
nor ( w8263 , w8262 , w7424 );
not ( w8264 , w8263 );
and ( w8265 , w8264 , w7428 );
not ( w8266 , w8265 );
and ( w8267 , w310 , w8266 );
and ( w8268 , w8267 , w8272 );
not ( w8269 , w8268 );
and ( w8270 , w8269 , w7428 );
nor ( w8271 , w310 , w8270 );
not ( w8272 , w7424 );
and ( w8273 , w8271 , w8272 );
not ( w8274 , w8273 );
and ( w8275 , w8274 , w7428 );
and ( w8276 , w8275 , w7458 );
and ( w8277 , w8276 , w7428 );
and ( w8278 , w8277 , w7458 );
and ( w8279 , w8278 , w7428 );
and ( w8280 , w8279 , w8275 );
not ( w8281 , w8280 );
and ( w8282 , w310 , w8281 );
not ( w8283 , w8282 );
and ( w8284 , w7445 , w8283 );
and ( w8285 , w8284 , w7459 );
and ( w8286 , w8285 , w7458 );
and ( w8287 , w8286 , w7428 );
and ( w8288 , w8287 , w20 );
nor ( w8289 , w8288 , w8074 );
and ( w8290 , w8289 , w12498 );
not ( w8291 , w8290 );
and ( w8292 , w8291 , w7459 );
and ( w8293 , w8292 , w8211 );
and ( w8294 , w8640 , w8293 );
and ( w8295 , w8294 , w11166 );
nor ( w8296 , w8295 , w19 );
not ( w8297 , w8296 );
and ( w8298 , w8297 , w8068 );
and ( w8299 , w8298 , w7458 );
and ( w8300 , w8299 , w7428 );
and ( w8301 , w8300 , w7418 );
and ( w8302 , w8301 , w7448 );
not ( w8303 , w8302 );
and ( w8304 , w8260 , w8303 );
not ( w8305 , w7513 );
and ( w8306 , w8304 , w8305 );
and ( w8307 , w8306 , w12144 );
and ( w8308 , w8307 , w12919 );
and ( w8309 , w8308 , w12142 );
and ( w8310 , w8309 , w8640 );
and ( w8311 , w8310 , w12921 );
nor ( w8312 , w7487 , w37 );
not ( w8313 , w8312 );
and ( w8314 , w8313 , w7459 );
nor ( w8315 , w8314 , w41 );
not ( w8316 , w8315 );
and ( w8317 , w8316 , w7459 );
nor ( w8318 , w8317 , w7522 );
not ( w8319 , w8318 );
and ( w8320 , w8319 , w7459 );
and ( w8321 , w8320 , w7810 );
and ( w8322 , w8321 , w7527 );
nor ( w8323 , w8322 , w20 );
and ( w8324 , w8323 , w485 );
and ( w8325 , w7522 , w12919 );
and ( w8326 , w12921 , w8325 );
not ( w8327 , w8326 );
and ( w8328 , w8327 , w485 );
not ( w8329 , w8328 );
and ( w8330 , w8329 , w7527 );
nor ( w8331 , w8330 , w8302 );
and ( w8332 , w8331 , w12921 );
and ( w8333 , w8332 , w11166 );
not ( w8334 , w8333 );
and ( w8335 , w8334 , w8109 );
and ( w8336 , w8335 , w8068 );
nor ( w8337 , w8336 , w7435 );
not ( w8338 , w8337 );
and ( w8339 , w8338 , w7428 );
and ( w8340 , w8339 , w7448 );
and ( w8341 , w8324 , w8408 );
and ( w8342 , w8341 , w11166 );
not ( w8343 , w8342 );
and ( w8344 , w8343 , w8109 );
nor ( w8345 , w8344 , w19 );
not ( w8346 , w8345 );
and ( w8347 , w8346 , w8068 );
and ( w8348 , w8347 , w7458 );
nor ( w8349 , w8348 , w7435 );
not ( w8350 , w8349 );
and ( w8351 , w8350 , w7428 );
and ( w8352 , w8351 , w7418 );
and ( w8353 , w8352 , w7448 );
not ( w8354 , w8311 );
and ( w8355 , w8354 , w8353 );
and ( w8356 , w8355 , w8109 );
and ( w8357 , w8356 , w12037 );
nor ( w8358 , w8083 , w31 );
not ( w8359 , w8358 );
and ( w8360 , w8359 , w7459 );
and ( w8361 , w8360 , w7504 );
and ( w8362 , w8361 , w7459 );
not ( w8363 , w35 );
and ( w8364 , w8362 , w8363 );
and ( w8365 , w8364 , w11347 );
nor ( w8366 , w8365 , w37 );
not ( w8367 , w8366 );
and ( w8368 , w8367 , w7459 );
and ( w8369 , w8368 , w11140 );
nor ( w8370 , w8369 , w41 );
nor ( w8371 , w8370 , w45 );
nor ( w8372 , w8193 , w8153 );
not ( w8373 , w8211 );
and ( w8374 , w8372 , w8373 );
and ( w8375 , w8374 , w8640 );
and ( w8376 , w8375 , w12921 );
and ( w8377 , w8376 , w11166 );
and ( w8378 , w8377 , w8848 );
not ( w8379 , w8378 );
and ( w8380 , w8379 , w8068 );
and ( w8381 , w8380 , w7458 );
and ( w8382 , w8381 , w7428 );
and ( w8383 , w8382 , w7418 );
and ( w8384 , w8383 , w7448 );
nor ( w8385 , w8371 , w8384 );
and ( w8386 , w8385 , w12144 );
and ( w8387 , w8386 , w12919 );
and ( w8388 , w8387 , w12142 );
not ( w8389 , w8388 );
and ( w8390 , w8389 , w7428 );
nor ( w8391 , w8390 , w485 );
and ( w8392 , w8391 , w12921 );
nor ( w8393 , w7487 , w37 );
not ( w8394 , w8393 );
and ( w8395 , w8394 , w7459 );
nor ( w8396 , w8395 , w41 );
not ( w8397 , w8396 );
and ( w8398 , w8397 , w7459 );
and ( w8399 , w8398 , w12117 );
and ( w8400 , w8399 , w7507 );
nor ( w8401 , w8400 , w7522 );
not ( w8402 , w8401 );
and ( w8403 , w8402 , w7810 );
and ( w8404 , w8403 , w7459 );
and ( w8405 , w8404 , w7527 );
not ( w8406 , w8405 );
and ( w8407 , w8406 , w485 );
not ( w8408 , w8340 );
and ( w8409 , w8407 , w8408 );
and ( w8410 , w8409 , w12921 );
and ( w8411 , w8410 , w11166 );
not ( w8412 , w8411 );
and ( w8413 , w8412 , w8109 );
nor ( w8414 , w8413 , w19 );
not ( w8415 , w8414 );
and ( w8416 , w8415 , w8068 );
and ( w8417 , w8416 , w7458 );
nor ( w8418 , w8417 , w7435 );
not ( w8419 , w8418 );
and ( w8420 , w8419 , w7428 );
and ( w8421 , w8420 , w7418 );
and ( w8422 , w8421 , w7448 );
not ( w8423 , w8392 );
and ( w8424 , w8423 , w8422 );
and ( w8425 , w8424 , w8109 );
and ( w8426 , w8425 , w12532 );
nor ( w8427 , w8426 , w19 );
not ( w8428 , w8427 );
and ( w8429 , w8428 , w8068 );
and ( w8430 , w8429 , w7458 );
nor ( w8431 , w8430 , w7435 );
not ( w8432 , w8431 );
and ( w8433 , w8432 , w7428 );
and ( w8434 , w8433 , w7418 );
and ( w8435 , w8434 , w7448 );
nor ( w8436 , w8357 , w8435 );
and ( w8437 , w8436 , w11166 );
not ( w8438 , w8437 );
and ( w8439 , w8438 , w8109 );
nor ( w8440 , w8439 , w19 );
not ( w8441 , w8440 );
and ( w8442 , w8441 , w8068 );
and ( w8443 , w8442 , w7458 );
and ( w8444 , w8443 , w7428 );
and ( w8445 , w8444 , w7418 );
and ( w8446 , w8445 , w7448 );
not ( w8447 , w8236 );
and ( w8448 , w8447 , w8446 );
nor ( w8449 , w8448 , w105 );
not ( w8450 , w8449 );
and ( w8451 , w8450 , w8109 );
nor ( w8452 , w8451 , w19 );
not ( w8453 , w8452 );
and ( w8454 , w8453 , w8068 );
and ( w8455 , w8454 , w7458 );
and ( w8456 , w8455 , w7428 );
and ( w8457 , w8456 , w7418 );
and ( w8458 , w8457 , w7448 );
not ( w8459 , w8222 );
and ( w8460 , w8459 , w8458 );
nor ( w8461 , w8460 , w105 );
and ( w8462 , w7401 , w8876 );
not ( w8463 , w8462 );
and ( w8464 , w8463 , w7448 );
not ( w8465 , w8461 );
and ( w8466 , w8465 , w8464 );
nor ( w8467 , w8466 , w19 );
not ( w8468 , w8467 );
and ( w8469 , w8468 , w8068 );
and ( w8470 , w8469 , w7458 );
nor ( w8471 , w8470 , w7435 );
not ( w8472 , w8471 );
and ( w8473 , w8472 , w7428 );
and ( w8474 , w8473 , w7418 );
and ( w8475 , w8474 , w7448 );
nor ( w8476 , w8217 , w8475 );
not ( w8477 , w8476 );
and ( w8478 , w8477 , w7459 );
nor ( w8479 , w8478 , w20 );
not ( w8480 , w8479 );
and ( w8481 , w8480 , w8458 );
nor ( w8482 , w8481 , w105 );
not ( w8483 , w8482 );
and ( w8484 , w8483 , w8464 );
nor ( w8485 , w8484 , w19 );
not ( w8486 , w8485 );
and ( w8487 , w8486 , w8068 );
and ( w8488 , w8487 , w7458 );
nor ( w8489 , w8488 , w7435 );
not ( w8490 , w8489 );
and ( w8491 , w8490 , w7428 );
and ( w8492 , w8491 , w7418 );
and ( w8493 , w8492 , w7448 );
and ( w8494 , w8081 , w8493 );
nor ( w8495 , w8494 , w105 );
not ( w8496 , w8495 );
and ( w8497 , w8496 , w8464 );
and ( w8498 , w8497 , w8109 );
nor ( w8499 , w8498 , w19 );
not ( w8500 , w8499 );
and ( w8501 , w8500 , w8068 );
and ( w8502 , w8501 , w7458 );
and ( w8503 , w8502 , w7428 );
and ( w8504 , w8503 , w7418 );
and ( w8505 , w8504 , w7448 );
not ( w8506 , w7789 );
and ( w8507 , w8506 , w8505 );
and ( w8508 , w8507 , w8493 );
and ( w8509 , w8508 , w8464 );
and ( w8510 , w8509 , w8109 );
nor ( w8511 , w8510 , w19 );
not ( w8512 , w8511 );
and ( w8513 , w8512 , w8068 );
and ( w8514 , w8513 , w7458 );
nor ( w8515 , w8514 , w7435 );
not ( w8516 , w8515 );
and ( w8517 , w8516 , w7428 );
and ( w8518 , w8517 , w7418 );
and ( w8519 , w8518 , w7448 );
and ( w8520 , w7781 , w8644 );
not ( w8521 , w8520 );
and ( w8522 , w8521 , w7458 );
nor ( w8523 , w8522 , w7435 );
not ( w8524 , w8523 );
and ( w8525 , w8524 , w7428 );
and ( w8526 , w8525 , w7448 );
not ( w8527 , w7780 );
and ( w8528 , w8527 , w8526 );
nor ( w8529 , w8528 , w48 );
not ( w8530 , w8529 );
and ( w8531 , w8530 , w7428 );
nor ( w8532 , w8531 , w20 );
and ( w8533 , w8532 , w8640 );
and ( w8534 , w8533 , w11166 );
and ( w8535 , w8534 , w8848 );
and ( w8536 , w7671 , w11140 );
nor ( w8537 , w8536 , w43 );
not ( w8538 , w8537 );
and ( w8539 , w8538 , w7592 );
and ( w8540 , w8539 , w12919 );
nor ( w8541 , w8540 , w48 );
nor ( w8542 , w18 , w20 );
not ( w8543 , w8542 );
and ( w8544 , w8543 , w384 );
not ( w8545 , w8544 );
and ( w8546 , w8545 , w7458 );
nor ( w8547 , w8546 , w7435 );
not ( w8548 , w8547 );
and ( w8549 , w8548 , w7428 );
and ( w8550 , w8549 , w7418 );
and ( w8551 , w8550 , w7448 );
not ( w8552 , w8541 );
and ( w8553 , w8552 , w8551 );
and ( w8554 , w8553 , w7459 );
and ( w8555 , w8554 , w7810 );
and ( w8556 , w8555 , w19 );
and ( w8557 , w8556 , w11166 );
not ( w8558 , w8557 );
and ( w8559 , w8558 , w19 );
and ( w8560 , w8559 , w8051 );
and ( w8561 , w8560 , w8634 );
not ( w8562 , w8561 );
and ( w8563 , w8562 , w8057 );
nor ( w8564 , w8563 , w8037 );
and ( w8565 , w8564 , w8594 );
and ( w8566 , w8565 , w8798 );
not ( w8567 , w8566 );
and ( w8568 , w8567 , w7459 );
not ( w8569 , w8568 );
and ( w8570 , w8569 , w255 );
nor ( w8571 , w7522 , w7513 );
and ( w8572 , w8571 , w12144 );
and ( w8573 , w8572 , w12142 );
not ( w8574 , w8573 );
and ( w8575 , w8574 , w7527 );
nor ( w8576 , w8575 , w20 );
and ( w8577 , w8576 , w485 );
nor ( w8578 , w7599 , w7452 );
nor ( w8579 , w8578 , w18 );
not ( w8580 , w8579 );
and ( w8581 , w8580 , w8526 );
nor ( w8582 , w8581 , w48 );
not ( w8583 , w8582 );
and ( w8584 , w8583 , w7428 );
nor ( w8585 , w8584 , w19 );
and ( w8586 , w8585 , w12921 );
and ( w8587 , w12921 , w7691 );
and ( w8588 , w8587 , w7597 );
and ( w8589 , w8588 , w12919 );
and ( w8590 , w8589 , w7940 );
and ( w8591 , w8590 , w7810 );
nor ( w8592 , w8591 , w8037 );
and ( w8593 , w19 , w8592 );
not ( w8594 , w5252 );
and ( w8595 , w8593 , w8594 );
and ( w8596 , w8595 , w8640 );
not ( w8597 , w8596 );
and ( w8598 , w8597 , w7459 );
and ( w8599 , w8598 , w7712 );
nor ( w8600 , w8599 , w8519 );
not ( w8601 , w8600 );
and ( w8602 , w8601 , w7458 );
and ( w8603 , w8602 , w7428 );
and ( w8604 , w8603 , w7418 );
and ( w8605 , w8604 , w7448 );
not ( w8606 , w8586 );
and ( w8607 , w8606 , w8605 );
nor ( w8608 , w8607 , w7449 );
and ( w8609 , w8608 , w8640 );
and ( w8610 , w8609 , w11166 );
not ( w8611 , w8610 );
and ( w8612 , w8611 , w7712 );
nor ( w8613 , w8612 , w8519 );
not ( w8614 , w8613 );
and ( w8615 , w8614 , w7458 );
nor ( w8616 , w8615 , w7435 );
not ( w8617 , w8616 );
and ( w8618 , w8617 , w7428 );
and ( w8619 , w8618 , w7418 );
and ( w8620 , w8619 , w7448 );
and ( w8621 , w8620 , w8605 );
nor ( w8622 , w8621 , w105 );
not ( w8623 , w8622 );
and ( w8624 , w8623 , w7712 );
nor ( w8625 , w8624 , w8519 );
not ( w8626 , w8625 );
and ( w8627 , w8626 , w7458 );
and ( w8628 , w8627 , w7428 );
and ( w8629 , w8628 , w7418 );
and ( w8630 , w8629 , w7448 );
not ( w8631 , w8577 );
and ( w8632 , w8631 , w8630 );
nor ( w8633 , w8632 , w19 );
not ( w8634 , w8060 );
and ( w8635 , w8634 , w105 );
not ( w8636 , w8037 );
and ( w8637 , w8635 , w8636 );
not ( w8638 , w8637 );
and ( w8639 , w8638 , w8630 );
not ( w8640 , w485 );
and ( w8641 , w8639 , w8640 );
nor ( w8642 , w8641 , w5252 );
and ( w8643 , w8642 , w8798 );
not ( w8644 , w8519 );
and ( w8645 , w8643 , w8644 );
not ( w8646 , w8645 );
and ( w8647 , w8646 , w7448 );
not ( w8648 , w8633 );
and ( w8649 , w8648 , w8647 );
nor ( w8650 , w8649 , w7549 );
not ( w8651 , w8650 );
and ( w8652 , w8651 , w7712 );
nor ( w8653 , w8652 , w8519 );
not ( w8654 , w8653 );
and ( w8655 , w8654 , w7458 );
nor ( w8656 , w8655 , w7435 );
not ( w8657 , w8656 );
and ( w8658 , w8657 , w7428 );
and ( w8659 , w8658 , w7418 );
and ( w8660 , w8659 , w7448 );
and ( w8661 , w8845 , w8660 );
nor ( w8662 , w8661 , w19 );
not ( w8663 , w8662 );
and ( w8664 , w8663 , w8647 );
nor ( w8665 , w8664 , w7549 );
not ( w8666 , w8665 );
and ( w8667 , w8666 , w7458 );
nor ( w8668 , w8667 , w7435 );
not ( w8669 , w8668 );
and ( w8670 , w8669 , w7428 );
and ( w8671 , w8670 , w7418 );
and ( w8672 , w8671 , w7448 );
not ( w8673 , w8570 );
and ( w8674 , w8673 , w8672 );
nor ( w8675 , w8674 , w8519 );
not ( w8676 , w8675 );
and ( w8677 , w8676 , w7458 );
nor ( w8678 , w8677 , w7435 );
not ( w8679 , w8678 );
and ( w8680 , w8679 , w7428 );
and ( w8681 , w8680 , w7418 );
and ( w8682 , w8681 , w7448 );
not ( w8683 , w8535 );
and ( w8684 , w8683 , w8682 );
nor ( w8685 , w8684 , w377 );
not ( w8686 , w8685 );
and ( w8687 , w8686 , w7459 );
not ( w8688 , w8687 );
and ( w8689 , w8688 , w255 );
not ( w8690 , w8689 );
and ( w8691 , w8690 , w8672 );
and ( w8692 , w8691 , w7712 );
nor ( w8693 , w8692 , w8519 );
not ( w8694 , w8693 );
and ( w8695 , w8694 , w7458 );
nor ( w8696 , w8695 , w7435 );
not ( w8697 , w8696 );
and ( w8698 , w8697 , w7428 );
and ( w8699 , w8698 , w7418 );
and ( w8700 , w8699 , w7448 );
not ( w8701 , w7779 );
and ( w8702 , w8701 , w8700 );
nor ( w8703 , w8702 , w19 );
not ( w8704 , w8703 );
and ( w8705 , w8704 , w8682 );
not ( w8706 , w8705 );
and ( w8707 , w8706 , w255 );
not ( w8708 , w8707 );
and ( w8709 , w8708 , w8672 );
nor ( w8710 , w8709 , w7746 );
not ( w8711 , w8710 );
and ( w8712 , w8711 , w7712 );
nor ( w8713 , w8712 , w8519 );
not ( w8714 , w8713 );
and ( w8715 , w8714 , w7458 );
nor ( w8716 , w8715 , w7435 );
not ( w8717 , w8716 );
and ( w8718 , w8717 , w7428 );
and ( w8719 , w8718 , w7418 );
and ( w8720 , w8719 , w7448 );
and ( w8721 , w8845 , w8720 );
nor ( w8722 , w8721 , w19 );
not ( w8723 , w8722 );
and ( w8724 , w8723 , w8682 );
not ( w8725 , w8724 );
and ( w8726 , w8725 , w255 );
not ( w8727 , w8726 );
and ( w8728 , w8727 , w8672 );
nor ( w8729 , w8728 , w7746 );
not ( w8730 , w8729 );
and ( w8731 , w8730 , w7712 );
nor ( w8732 , w8731 , w8519 );
not ( w8733 , w8732 );
and ( w8734 , w8733 , w7458 );
nor ( w8735 , w8734 , w7435 );
not ( w8736 , w8735 );
and ( w8737 , w8736 , w7428 );
and ( w8738 , w8737 , w7418 );
and ( w8739 , w8738 , w7448 );
not ( w8740 , w8739 );
and ( w8741 , w7771 , w8740 );
not ( w8742 , w8741 );
and ( w8743 , w8742 , w7458 );
nor ( w8744 , w8743 , w7435 );
not ( w8745 , w8744 );
and ( w8746 , w8745 , w7428 );
and ( w8747 , w8746 , w7418 );
and ( w8748 , w8747 , w7448 );
not ( w8749 , w7764 );
and ( w8750 , w8749 , w8748 );
nor ( w8751 , w8750 , w8739 );
not ( w8752 , w8751 );
and ( w8753 , w8752 , w7458 );
nor ( w8754 , w8753 , w7435 );
not ( w8755 , w8754 );
and ( w8756 , w8755 , w7428 );
and ( w8757 , w8756 , w7418 );
and ( w8758 , w8757 , w7448 );
nor ( w8759 , w7713 , w8758 );
not ( w8760 , w8759 );
and ( w8761 , w8760 , w7458 );
nor ( w8762 , w8761 , w7435 );
not ( w8763 , w8762 );
and ( w8764 , w8763 , w7428 );
and ( w8765 , w8764 , w7418 );
and ( w8766 , w8765 , w7448 );
and ( w8767 , w7608 , w8766 );
nor ( w8768 , w8767 , w20 );
and ( w8769 , w8768 , w12142 );
not ( w8770 , w8769 );
and ( w8771 , w8770 , w7428 );
and ( w8772 , w8771 , w11166 );
nor ( w8773 , w8772 , w7449 );
nor ( w8774 , w8773 , w485 );
nor ( w8775 , w8774 , w8758 );
not ( w8776 , w8775 );
and ( w8777 , w8776 , w7458 );
nor ( w8778 , w8777 , w7435 );
not ( w8779 , w8778 );
and ( w8780 , w8779 , w7428 );
and ( w8781 , w8780 , w7448 );
and ( w8782 , w7597 , w8781 );
and ( w8783 , w310 , w7585 );
not ( w8784 , w8783 );
and ( w8785 , w8784 , w20 );
not ( w8786 , w8785 );
and ( w8787 , w8786 , w7458 );
nor ( w8788 , w8787 , w7435 );
not ( w8789 , w8788 );
and ( w8790 , w8789 , w7428 );
and ( w8791 , w8790 , w7448 );
and ( w8792 , w8782 , w8791 );
and ( w8793 , w8792 , w19 );
and ( w8794 , w8793 , w377 );
and ( w8795 , w8794 , w11166 );
nor ( w8796 , w8795 , w7449 );
and ( w8797 , w8796 , w7761 );
not ( w8798 , w7760 );
and ( w8799 , w8797 , w8798 );
not ( w8800 , w8799 );
and ( w8801 , w8800 , w7459 );
and ( w8802 , w8801 , w7712 );
nor ( w8803 , w8802 , w8758 );
not ( w8804 , w8803 );
and ( w8805 , w8804 , w7458 );
nor ( w8806 , w8805 , w7435 );
not ( w8807 , w8806 );
and ( w8808 , w8807 , w7428 );
and ( w8809 , w8808 , w7418 );
and ( w8810 , w8809 , w7448 );
not ( w8811 , w7557 );
and ( w8812 , w8811 , w8810 );
nor ( w8813 , w8812 , w7746 );
not ( w8814 , w8813 );
and ( w8815 , w8814 , w7712 );
nor ( w8816 , w8815 , w8758 );
not ( w8817 , w8816 );
and ( w8818 , w8817 , w7458 );
nor ( w8819 , w8818 , w7435 );
not ( w8820 , w8819 );
and ( w8821 , w8820 , w7428 );
and ( w8822 , w8821 , w7418 );
and ( w8823 , w8822 , w7448 );
nor ( w8824 , w8823 , w7449 );
and ( w8825 , w8824 , w12142 );
not ( w8826 , w8825 );
and ( w8827 , w8826 , w7428 );
nor ( w8828 , w8827 , w20 );
not ( w8829 , w7555 );
and ( w8830 , w8828 , w8829 );
and ( w8831 , w8830 , w8848 );
not ( w8832 , w8831 );
and ( w8833 , w8832 , w8810 );
nor ( w8834 , w8833 , w7746 );
not ( w8835 , w8834 );
and ( w8836 , w8835 , w7712 );
nor ( w8837 , w8836 , w8758 );
not ( w8838 , w8837 );
and ( w8839 , w8838 , w7458 );
nor ( w8840 , w8839 , w7435 );
not ( w8841 , w8840 );
and ( w8842 , w8841 , w7428 );
and ( w8843 , w8842 , w7418 );
and ( w8844 , w8843 , w7448 );
not ( w8845 , w7401 );
and ( w8846 , w8845 , w8844 );
nor ( w8847 , w8846 , w7549 );
not ( w8848 , w19 );
and ( w8849 , w8847 , w8848 );
not ( w8850 , w8849 );
and ( w8851 , w8850 , w8810 );
and ( w8852 , w8851 , w7458 );
nor ( w8853 , w8852 , w7435 );
not ( w8854 , w8853 );
and ( w8855 , w8854 , w7428 );
and ( w8856 , w8855 , w7418 );
and ( w8857 , w8856 , w7448 );
and ( w8858 , w12080 , w8857 );
nor ( w8859 , w8858 , w8758 );
not ( w8860 , w8859 );
and ( w8861 , w8860 , w7448 );
nor ( w8862 , w8861 , w7435 );
not ( w8863 , w8862 );
and ( w8864 , w8863 , w7448 );
nor ( w8865 , w8861 , w8864 );
and ( w8866 , w7445 , w7458 );
not ( w8867 , w7455 );
and ( w8868 , g6 , w8867 );
nor ( w8869 , w8868 , g5 );
nor ( w8870 , g7 , w8869 );
not ( w8871 , w8870 );
and ( w8872 , w8871 , w8865 );
nor ( w8873 , w8872 , g5 );
not ( w8874 , w8873 );
and ( w8875 , w8874 , w8865 );
not ( w8876 , w7435 );
and ( w8877 , w8875 , w8876 );
not ( w8878 , w8877 );
and ( w8879 , w8878 , w7428 );
and ( w8880 , w8866 , w8879 );
not ( w8881 , w52 );
and ( w8882 , w8880 , w8881 );
and ( w8883 , w7448 , w8879 );
nor ( w8884 , w8882 , w8883 );
not ( w8885 , w8884 );
and ( w8886 , w8885 , w8880 );
and ( w8887 , w8886 , w8879 );
and ( w8888 , w8887 , w8880 );
and ( w8889 , w8888 , w8879 );
and ( w8890 , w8889 , w8880 );
and ( w8891 , w8890 , w8879 );
and ( w8892 , w8891 , w13331 );
and ( w8893 , w8892 , w13333 );
and ( w8894 , w8891 , w13204 );
and ( w8895 , w8894 , w13206 );
and ( w8896 , w8895 , w8891 );
and ( w8897 , w8896 , w13204 );
and ( w8898 , w8897 , w13206 );
and ( w8899 , w8893 , w8898 );
and ( w8900 , w8890 , g48 );
and ( w8901 , w8900 , w13206 );
and ( w8902 , w8890 , w13204 );
and ( w8903 , w8902 , g31 );
and ( w8904 , w8903 , w8890 );
and ( w8905 , w8904 , w13204 );
nor ( w8906 , w8901 , w8905 );
and ( w8907 , w10949 , w8890 );
and ( w8908 , w8891 , g48 );
and ( w8909 , w8908 , g31 );
nor ( w8910 , w8907 , w8909 );
and ( w8911 , w9761 , w8891 );
and ( w8912 , w8894 , g31 );
nor ( w8913 , w8908 , w8912 );
and ( w8914 , w8911 , w10955 );
and ( w8915 , w8914 , w8891 );
and ( w8916 , w8915 , w8890 );
and ( w8917 , w8916 , w8891 );
and ( w8918 , w8917 , w8879 );
and ( w8919 , w8879 , w11795 );
and ( w8920 , w8919 , w11797 );
not ( w8921 , w8883 );
and ( w8922 , w8921 , w8865 );
and ( w8923 , w9601 , w8922 );
and ( w8924 , w8918 , w10662 );
and ( w8925 , w8879 , w9195 );
and ( w8926 , w8925 , w9197 );
not ( w8927 , w8926 );
and ( w8928 , w8927 , w8922 );
and ( w8929 , w8928 , w8865 );
and ( w8930 , w8879 , w9354 );
and ( w8931 , w8930 , w9356 );
not ( w8932 , w8931 );
and ( w8933 , w8932 , w8865 );
and ( w8934 , w8929 , w8933 );
and ( w8935 , w8891 , w9380 );
and ( w8936 , w8935 , w13321 );
and ( w8937 , w8934 , w10994 );
and ( w8938 , w8879 , w9053 );
and ( w8939 , w8938 , w9049 );
not ( w8940 , w8939 );
and ( w8941 , w8940 , w8922 );
and ( w8942 , w8922 , g41 );
and ( w8943 , w8942 , g15 );
not ( w8944 , w8943 );
and ( w8945 , w8944 , w8891 );
and ( w8946 , w8945 , w9053 );
not ( w8947 , w8946 );
and ( w8948 , w8947 , w8865 );
and ( w8949 , w8948 , g17 );
and ( w8950 , w8942 , g40 );
and ( w8951 , w8950 , g15 );
not ( w8952 , w8951 );
and ( w8953 , w8952 , w8891 );
not ( w8954 , w8949 );
and ( w8955 , w8954 , w8953 );
not ( w8956 , w8955 );
and ( w8957 , w8956 , w8922 );
and ( w8958 , w8891 , w10969 );
and ( w8959 , w8958 , w8879 );
and ( w8960 , w8959 , w8891 );
and ( w8961 , w8960 , g40 );
and ( w8962 , w8961 , w9049 );
not ( w8963 , w8962 );
and ( w8964 , w8963 , w8922 );
and ( w8965 , w8959 , w9053 );
and ( w8966 , w8965 , g17 );
not ( w8967 , w8966 );
and ( w8968 , w8967 , w8922 );
and ( w8969 , w8964 , w8968 );
and ( w8970 , w8941 , w8969 );
and ( w8971 , w8922 , w8970 );
not ( w8972 , w8971 );
and ( w8973 , w8972 , w8891 );
and ( w8974 , w8865 , g37 );
and ( w8975 , w8974 , g19 );
not ( w8976 , w8975 );
and ( w8977 , w8976 , w8891 );
and ( w8978 , w8973 , w8977 );
and ( w8979 , w8937 , w10852 );
not ( w8980 , w8979 );
and ( w8981 , w8980 , w8879 );
and ( w8982 , w8981 , w8891 );
and ( w8983 , g38 , g25 );
not ( w8984 , w8983 );
and ( w8985 , w8984 , w8891 );
not ( w8986 , g44 );
and ( w8987 , w8879 , w8986 );
and ( w8988 , w8987 , w13050 );
nor ( w8989 , w8985 , w8988 );
and ( w8990 , w8982 , w10999 );
not ( w8991 , w8990 );
and ( w8992 , w8991 , w8865 );
and ( w8993 , w8879 , w12962 );
and ( w8994 , w8993 , w12964 );
and ( w8995 , w8992 , w10276 );
not ( w8996 , w8987 );
and ( w8997 , w8996 , g27 );
nor ( w8998 , w8995 , w8997 );
not ( w8999 , w8998 );
and ( w9000 , w8999 , w8865 );
and ( w9001 , w9000 , w8922 );
and ( w9002 , w10568 , w8922 );
and ( w9003 , w9001 , w9002 );
and ( w9004 , w8865 , g46 );
not ( w9005 , w9004 );
and ( w9006 , w9005 , w8879 );
not ( w9007 , w9006 );
and ( w9008 , w9007 , g9 );
nor ( w9009 , w9003 , w9008 );
not ( w9010 , g46 );
and ( w9011 , w8879 , w9010 );
and ( w9012 , w9011 , w13590 );
and ( w9013 , w11004 , w8922 );
nor ( w9014 , w9008 , w9013 );
not ( w9015 , w9014 );
and ( w9016 , w9015 , w8922 );
not ( w9017 , w9009 );
and ( w9018 , w9017 , w9016 );
not ( w9019 , w8919 );
and ( w9020 , w9019 , g13 );
and ( w9021 , w8923 , w9020 );
nor ( w9022 , w9018 , w9021 );
not ( w9023 , w9022 );
and ( w9024 , w9023 , w8865 );
and ( w9025 , w9024 , w8922 );
and ( w9026 , w8879 , w13474 );
and ( w9027 , w9026 , w13477 );
and ( w9028 , w10905 , w8922 );
nor ( w9029 , w9025 , w9028 );
and ( w9030 , w8922 , g39 );
not ( w9031 , w9030 );
and ( w9032 , w9031 , w8879 );
not ( w9033 , w9032 );
and ( w9034 , w9033 , g13 );
and ( w9035 , w9034 , w9020 );
and ( w9036 , w8928 , w8933 );
and ( w9037 , w8977 , w10510 );
not ( w9038 , w9037 );
and ( w9039 , w9038 , w8922 );
and ( w9040 , w9036 , w9039 );
nor ( w9041 , w9040 , w8989 );
and ( w9042 , w9041 , w8891 );
and ( w9043 , w9042 , w10949 );
and ( w9044 , w8890 , w9053 );
and ( w9045 , w9044 , w9049 );
not ( w9046 , w9045 );
and ( w9047 , w9046 , w8922 );
and ( w9048 , w8958 , g40 );
not ( w9049 , g17 );
and ( w9050 , w9048 , w9049 );
not ( w9051 , w9050 );
and ( w9052 , w9051 , w8922 );
not ( w9053 , g40 );
and ( w9054 , w8958 , w9053 );
and ( w9055 , w9054 , g17 );
not ( w9056 , w9055 );
and ( w9057 , w9056 , w8922 );
and ( w9058 , w9052 , w9057 );
and ( w9059 , w9047 , w9058 );
and ( w9060 , w8891 , w10508 );
and ( w9061 , w9060 , w10510 );
not ( w9062 , w9039 );
and ( w9063 , w9061 , w9062 );
not ( w9064 , w9063 );
and ( w9065 , w9064 , w8922 );
and ( w9066 , w8891 , w9354 );
and ( w9067 , w9066 , w9356 );
not ( w9068 , w9067 );
and ( w9069 , w9068 , w8865 );
and ( w9070 , w9065 , w9069 );
not ( w9071 , w9070 );
and ( w9072 , w9071 , w8891 );
not ( w9073 , w9072 );
and ( w9074 , w9073 , w8928 );
not ( w9075 , w9074 );
and ( w9076 , w9075 , w8891 );
and ( w9077 , w9043 , w9076 );
not ( w9078 , w9077 );
and ( w9079 , w9078 , w8922 );
not ( w9080 , w9079 );
and ( w9081 , w9080 , w8891 );
not ( w9082 , w9081 );
and ( w9083 , w9082 , w8865 );
nor ( w9084 , g43 , g23 );
and ( w9085 , w11732 , w8891 );
not ( w9086 , w9083 );
and ( w9087 , w9086 , w9085 );
not ( w9088 , w9087 );
and ( w9089 , w9088 , w8922 );
not ( w9090 , w9089 );
and ( w9091 , w9090 , w8891 );
not ( w9092 , w9091 );
and ( w9093 , w9092 , w8865 );
not ( w9094 , w9093 );
and ( w9095 , w9094 , w8891 );
and ( w9096 , w9095 , w8985 );
and ( w9097 , w9096 , w8891 );
not ( w9098 , w9097 );
and ( w9099 , w9098 , w8865 );
nor ( w9100 , w9099 , w8997 );
not ( w9101 , w9100 );
and ( w9102 , w9101 , w8922 );
and ( w9103 , w9102 , w8865 );
and ( w9104 , w9103 , w8922 );
and ( w9105 , w9104 , w9002 );
not ( w9106 , w9105 );
and ( w9107 , w9106 , w8891 );
nor ( w9108 , g44 , g27 );
and ( w9109 , w13528 , w8891 );
and ( w9110 , w9107 , w9109 );
and ( w9111 , w9110 , w8891 );
and ( w9112 , w9111 , w8879 );
and ( w9113 , w13045 , w8891 );
and ( w9114 , w9112 , w9113 );
not ( w9115 , w9114 );
and ( w9116 , w9115 , w8922 );
not ( w9117 , w9116 );
and ( w9118 , w9117 , w8891 );
and ( w9119 , w8922 , w13474 );
and ( w9120 , w9119 , w13477 );
not ( w9121 , w9120 );
and ( w9122 , w9121 , w8879 );
and ( w9123 , w9118 , w9122 );
and ( w9124 , w8879 , w11217 );
and ( w9125 , w9124 , w13211 );
and ( w9126 , w9758 , w8922 );
not ( w9127 , w9123 );
and ( w9128 , w9127 , w9126 );
and ( w9129 , g47 , w8879 );
nor ( w9130 , w9129 , g33 );
not ( w9131 , w9124 );
and ( w9132 , w9131 , g33 );
nor ( w9133 , w9130 , w9132 );
not ( w9134 , w9128 );
and ( w9135 , w9134 , w9133 );
and ( w9136 , w10276 , w8865 );
nor ( w9137 , w9136 , w8997 );
not ( w9138 , w9137 );
and ( w9139 , w9138 , w8865 );
and ( w9140 , w9139 , w8922 );
and ( w9141 , w9140 , w9002 );
nor ( w9142 , w9141 , w9008 );
not ( w9143 , w9142 );
and ( w9144 , w9143 , w8922 );
and ( w9145 , w9144 , w8923 );
and ( w9146 , w9145 , w9016 );
nor ( w9147 , w9146 , w9021 );
not ( w9148 , w9147 );
and ( w9149 , w9148 , w8865 );
and ( w9150 , w9149 , w8922 );
nor ( w9151 , w9150 , w9028 );
not ( w9152 , w8897 );
and ( w9153 , w9152 , w8922 );
and ( w9154 , w9153 , w10329 );
and ( w9155 , w9154 , w8922 );
not ( w9156 , w9155 );
and ( w9157 , w9156 , w8893 );
and ( w9158 , w8928 , w8970 );
and ( w9159 , w9141 , w10414 );
not ( w9160 , w9159 );
and ( w9161 , w9160 , w8891 );
not ( w9162 , w9008 );
and ( w9163 , w9161 , w9162 );
nor ( w9164 , w9163 , w8936 );
not ( w9165 , w9164 );
and ( w9166 , w9165 , w8879 );
and ( w9167 , w9166 , w8891 );
not ( w9168 , w9167 );
and ( w9169 , w9168 , w8922 );
and ( w9170 , w9169 , w8923 );
and ( w9171 , w9170 , w9016 );
and ( w9172 , w9136 , w8989 );
nor ( w9173 , w9172 , w8997 );
not ( w9174 , w9173 );
and ( w9175 , w9174 , w8865 );
and ( w9176 , w9175 , w8922 );
and ( w9177 , w9176 , w9002 );
nor ( w9178 , w9177 , w9008 );
and ( w9179 , w10680 , w9016 );
and ( w9180 , w9179 , w8865 );
not ( w9181 , w9180 );
and ( w9182 , w9181 , w9027 );
nor ( w9183 , w8989 , w8997 );
nor ( w9184 , w9183 , w9012 );
not ( w9185 , w9184 );
and ( w9186 , w9185 , w8891 );
not ( w9187 , w9011 );
and ( w9188 , w9187 , g9 );
nor ( w9189 , w9184 , w9188 );
not ( w9190 , w9189 );
and ( w9191 , w8923 , w9190 );
and ( w9192 , w8879 , g36 );
and ( w9193 , w9192 , g11 );
and ( w9194 , w9191 , w10615 );
not ( w9195 , g37 );
and ( w9196 , w8891 , w9195 );
not ( w9197 , g19 );
and ( w9198 , w9196 , w9197 );
and ( w9199 , w8922 , w10987 );
and ( w9200 , w9199 , w8957 );
not ( w9201 , w9200 );
and ( w9202 , w9201 , w8977 );
and ( w9203 , w9202 , w8891 );
not ( w9204 , w8930 );
and ( w9205 , w9204 , g21 );
and ( w9206 , w9203 , w10200 );
not ( w9207 , w9206 );
and ( w9208 , w9207 , w8865 );
and ( w9209 , w9208 , w9069 );
and ( w9210 , w9209 , w10994 );
not ( w9211 , w9210 );
and ( w9212 , w9211 , w8985 );
and ( w9213 , g43 , g23 );
and ( w9214 , w13492 , w8891 );
and ( w9215 , w9212 , w9214 );
and ( w9216 , w8891 , w8994 );
nor ( w9217 , w9216 , w8988 );
not ( w9218 , w9217 );
and ( w9219 , w9218 , w8891 );
nor ( w9220 , w9215 , w9219 );
and ( w9221 , w9219 , w10978 );
nor ( w9222 , w9221 , w8988 );
not ( w9223 , w9222 );
and ( w9224 , w9223 , w8891 );
and ( w9225 , w9220 , w9431 );
not ( w9226 , w9225 );
and ( w9227 , w9226 , w8891 );
and ( w9228 , w9227 , w10978 );
and ( w9229 , w9228 , w9113 );
nor ( w9230 , w9229 , w9012 );
not ( w9231 , w9230 );
and ( w9232 , w9231 , w8891 );
nor ( w9233 , w9232 , w9133 );
not ( w9234 , w9233 );
and ( w9235 , w9234 , w8891 );
and ( w9236 , g45 , w8879 );
nor ( w9237 , w9236 , g29 );
and ( w9238 , w9235 , w10188 );
nor ( w9239 , w9238 , w9027 );
not ( w9240 , w9026 );
and ( w9241 , w9240 , g11 );
and ( w9242 , w9239 , w9241 );
not ( w9243 , w9242 );
and ( w9244 , w9243 , w8891 );
not ( w9245 , w9194 );
and ( w9246 , w9245 , w9244 );
nor ( w9247 , w9246 , w9133 );
and ( w9248 , w8879 , g39 );
and ( w9249 , w9248 , g13 );
and ( w9250 , w9247 , w11022 );
not ( w9251 , w9250 );
and ( w9252 , w9251 , w8891 );
not ( w9253 , w8993 );
and ( w9254 , w9253 , g25 );
not ( w9255 , w9254 );
and ( w9256 , w9255 , w8879 );
and ( w9257 , w9256 , w8891 );
and ( w9258 , w9257 , w8936 );
nor ( w9259 , w9258 , w8994 );
nor ( w9260 , w9259 , w8997 );
nor ( w9261 , w8988 , w9260 );
and ( w9262 , w8891 , w9198 );
not ( w9263 , w9262 );
and ( w9264 , w9263 , w8865 );
and ( w9265 , w9264 , w8933 );
not ( w9266 , w9265 );
and ( w9267 , w9266 , w8891 );
and ( w9268 , w9267 , w10200 );
and ( w9269 , w9268 , w9214 );
nor ( w9270 , w9269 , w8936 );
not ( w9271 , w9270 );
and ( w9272 , w9271 , w8879 );
and ( w9273 , w9272 , w8891 );
and ( w9274 , w9273 , w9252 );
not ( w9275 , w9274 );
and ( w9276 , w9261 , w9275 );
and ( w9277 , w9276 , w11004 );
not ( w9278 , w9277 );
and ( w9279 , w9278 , w8891 );
and ( w9280 , w9279 , w8879 );
and ( w9281 , w9280 , w9113 );
nor ( w9282 , w9281 , w9193 );
not ( w9283 , w9282 );
and ( w9284 , w9283 , w9244 );
and ( w9285 , w9129 , g33 );
nor ( w9286 , w9125 , w9285 );
and ( w9287 , w9284 , w10234 );
nor ( w9288 , w9287 , w9249 );
not ( w9289 , w9288 );
and ( w9290 , w9289 , w8891 );
nor ( w9291 , w9252 , w9290 );
nor ( w9292 , w9291 , w9286 );
and ( w9293 , w9186 , w9292 );
nor ( w9294 , w9293 , w8988 );
nor ( w9295 , w9294 , w9188 );
nor ( w9296 , w9295 , w9193 );
not ( w9297 , w9296 );
and ( w9298 , w9297 , w9244 );
nor ( w9299 , w9298 , w9249 );
not ( w9300 , w9299 );
and ( w9301 , w9300 , w8891 );
and ( w9302 , w9301 , w10188 );
and ( w9303 , w9302 , w10234 );
nor ( w9304 , w9182 , w9303 );
and ( w9305 , w9304 , w8922 );
and ( w9306 , w9305 , w8923 );
and ( w9307 , w9306 , w8865 );
not ( w9308 , w9307 );
and ( w9309 , w9308 , w9244 );
nor ( w9310 , w9309 , w9249 );
not ( w9311 , w9310 );
and ( w9312 , w9311 , w8891 );
and ( w9313 , w9312 , w10234 );
not ( w9314 , w9171 );
and ( w9315 , w9314 , w9313 );
not ( w9316 , w9315 );
and ( w9317 , w9316 , w8865 );
and ( w9318 , w9317 , w8922 );
nor ( w9319 , w9318 , w9241 );
nor ( w9320 , w9319 , w9122 );
not ( w9321 , w9320 );
and ( w9322 , w9321 , w9027 );
nor ( w9323 , w9262 , w9260 );
and ( w9324 , w9323 , w8922 );
and ( w9325 , w9324 , w8970 );
not ( w9326 , w9260 );
and ( w9327 , w8865 , w9326 );
and ( w9328 , w9327 , w10414 );
not ( w9329 , w9328 );
and ( w9330 , w9329 , w8891 );
and ( w9331 , w9330 , w9303 );
and ( w9332 , w9331 , w10200 );
nor ( w9333 , w9332 , w9012 );
not ( w9334 , w9333 );
and ( w9335 , w9334 , w8891 );
and ( w9336 , w9335 , w9122 );
nor ( w9337 , w9336 , w8988 );
nor ( w9338 , w9337 , w9188 );
not ( w9339 , w9338 );
and ( w9340 , w9339 , w8922 );
and ( w9341 , w9340 , w8923 );
and ( w9342 , w9341 , w10615 );
not ( w9343 , w9342 );
and ( w9344 , w9343 , w9244 );
and ( w9345 , w9344 , w8891 );
and ( w9346 , w9345 , w10179 );
not ( w9347 , w9346 );
and ( w9348 , w9347 , w8922 );
and ( w9349 , w9348 , w8865 );
and ( w9350 , w9349 , w8933 );
and ( w9351 , w10130 , w9313 );
not ( w9352 , w9351 );
and ( w9353 , w9352 , w8865 );
not ( w9354 , g42 );
and ( w9355 , w9353 , w9354 );
not ( w9356 , g21 );
and ( w9357 , w9355 , w9356 );
not ( w9358 , w9357 );
and ( w9359 , w9358 , w8879 );
and ( w9360 , w9359 , w8891 );
and ( w9361 , w8865 , w9205 );
not ( w9362 , w9361 );
and ( w9363 , w9362 , w8879 );
and ( w9364 , w9363 , w9380 );
not ( w9365 , w9364 );
and ( w9366 , w9365 , w8865 );
and ( w9367 , w9366 , g23 );
and ( w9368 , w8922 , w9205 );
not ( w9369 , w9368 );
and ( w9370 , w9369 , w8891 );
nor ( w9371 , w9370 , g23 );
not ( w9372 , w9371 );
and ( w9373 , w9372 , w8891 );
not ( w9374 , w9367 );
and ( w9375 , w9374 , w9373 );
not ( w9376 , w9375 );
and ( w9377 , w9376 , g23 );
not ( w9378 , w9377 );
and ( w9379 , w9378 , w8891 );
not ( w9380 , g43 );
and ( w9381 , w8879 , w9380 );
and ( w9382 , w9381 , w13321 );
not ( w9383 , w9382 );
and ( w9384 , w9383 , w8922 );
and ( w9385 , w9384 , g42 );
not ( w9386 , w9385 );
and ( w9387 , w9386 , w8879 );
not ( w9388 , w9387 );
and ( w9389 , w9388 , g21 );
not ( w9390 , w9389 );
and ( w9391 , w9390 , w8891 );
and ( w9392 , w9391 , w8879 );
and ( w9393 , w9392 , w12962 );
and ( w9394 , w9393 , w8891 );
and ( w9395 , w9394 , w9214 );
not ( w9396 , w9395 );
and ( w9397 , w9396 , w8922 );
and ( w9398 , w9397 , g25 );
and ( w9399 , w9391 , w9214 );
not ( w9400 , w9399 );
and ( w9401 , w9400 , w8922 );
and ( w9402 , w9401 , g38 );
not ( w9403 , w9402 );
and ( w9404 , w9403 , w8879 );
not ( w9405 , w9398 );
and ( w9406 , w9405 , w9404 );
not ( w9407 , w9406 );
and ( w9408 , w9407 , w8922 );
nor ( w9409 , w9408 , w8997 );
not ( w9410 , w9409 );
and ( w9411 , w9410 , w8865 );
and ( w9412 , w9411 , w8922 );
and ( w9413 , w9412 , w9002 );
nor ( w9414 , w9413 , w9008 );
not ( w9415 , w9414 );
and ( w9416 , w9415 , w9016 );
and ( w9417 , w9416 , w8865 );
and ( w9418 , w9417 , w13474 );
and ( w9419 , w9418 , w13477 );
not ( w9420 , w9419 );
and ( w9421 , w9420 , w8879 );
and ( w9422 , w8891 , w10978 );
and ( w9423 , w9422 , w8879 );
and ( w9424 , w8985 , w8936 );
not ( w9425 , w9424 );
and ( w9426 , w9425 , w9205 );
not ( w9427 , w9426 );
and ( w9428 , w9427 , w8891 );
and ( w9429 , w9428 , w9214 );
nor ( w9430 , w9429 , w9219 );
not ( w9431 , w9224 );
and ( w9432 , w9430 , w9431 );
not ( w9433 , w9432 );
and ( w9434 , w9433 , w8891 );
and ( w9435 , w9434 , w10978 );
and ( w9436 , w9435 , w9113 );
nor ( w9437 , w9436 , w9012 );
not ( w9438 , w9437 );
and ( w9439 , w9438 , w8891 );
and ( w9440 , w9423 , w9439 );
and ( w9441 , w9440 , w9113 );
nor ( w9442 , w9441 , w9012 );
not ( w9443 , w9442 );
and ( w9444 , w9443 , w8891 );
nor ( w9445 , w9444 , w9193 );
nor ( w9446 , w8895 , w8909 );
not ( w9447 , w9446 );
and ( w9448 , w9447 , w9439 );
and ( w9449 , w9448 , w8893 );
not ( w9450 , w9449 );
and ( w9451 , w9450 , w9241 );
not ( w9452 , w9451 );
and ( w9453 , w9452 , w8891 );
not ( w9454 , w9445 );
and ( w9455 , w9454 , w9453 );
and ( w9456 , w9455 , w8879 );
and ( w9457 , w9456 , w8891 );
nor ( w9458 , w9248 , g13 );
and ( w9459 , w9457 , w11029 );
nor ( w9460 , w9459 , w9249 );
not ( w9461 , w9460 );
and ( w9462 , w9461 , w8891 );
and ( w9463 , w9462 , w8893 );
and ( w9464 , w8891 , w9435 );
and ( w9465 , w9464 , w10978 );
nor ( w9466 , w9465 , w9012 );
not ( w9467 , w9466 );
and ( w9468 , w9467 , w8879 );
and ( w9469 , w9468 , w8891 );
and ( w9470 , w9469 , w8879 );
and ( w9471 , w9470 , w9113 );
nor ( w9472 , w8920 , w9471 );
nor ( w9473 , w9472 , w9241 );
and ( w9474 , w9473 , w10179 );
and ( w9475 , w8920 , w9499 );
and ( w9476 , w9471 , w10179 );
and ( w9477 , w9476 , w9499 );
nor ( w9478 , w9477 , w9027 );
not ( w9479 , w9475 );
and ( w9480 , w9479 , w9478 );
and ( w9481 , w9464 , w8879 );
and ( w9482 , w9481 , w8891 );
and ( w9483 , w9482 , w10978 );
and ( w9484 , w8891 , w9483 );
and ( w9485 , w9484 , w8879 );
nor ( w9486 , w9485 , w9471 );
not ( w9487 , w9486 );
and ( w9488 , w9487 , w9113 );
not ( w9489 , w9488 );
and ( w9490 , w9489 , w9478 );
and ( w9491 , w8891 , w10955 );
and ( w9492 , w10200 , w8891 );
and ( w9493 , w9492 , w9214 );
nor ( w9494 , w9493 , w8988 );
not ( w9495 , w9494 );
and ( w9496 , w9495 , w8891 );
and ( w9497 , w9496 , w8879 );
and ( w9498 , w9497 , w9113 );
not ( w9499 , w9241 );
and ( w9500 , w9498 , w9499 );
nor ( w9501 , w9500 , w9439 );
and ( w9502 , w9501 , w11004 );
not ( w9503 , w9502 );
and ( w9504 , w9503 , w8891 );
nor ( w9505 , w9504 , w9027 );
not ( w9506 , w9505 );
and ( w9507 , w9491 , w9506 );
and ( w9508 , w9507 , w8879 );
and ( w9509 , w9508 , w8891 );
and ( w9510 , w9509 , w11029 );
and ( w9511 , w9510 , w8891 );
nor ( w9512 , w9511 , w9285 );
and ( w9513 , w9512 , w9758 );
and ( w9514 , w8891 , w11795 );
and ( w9515 , w9514 , w11797 );
and ( w9516 , w9515 , w8891 );
and ( w9517 , w9516 , w10179 );
nor ( w9518 , w9012 , w9260 );
and ( w9519 , w9518 , w10568 );
nor ( w9520 , w9519 , w9188 );
and ( w9521 , w8988 , w9551 );
nor ( w9522 , w9520 , w9521 );
and ( w9523 , w9601 , w9522 );
nor ( w9524 , w9523 , w9020 );
nor ( w9525 , w9524 , w9193 );
and ( w9526 , w9525 , w9205 );
not ( w9527 , w9526 );
and ( w9528 , w9527 , w8891 );
and ( w9529 , w9528 , w9214 );
nor ( w9530 , w9260 , w8994 );
nor ( w9531 , w9530 , w8997 );
nor ( w9532 , w9529 , w9531 );
and ( w9533 , w9532 , w10568 );
and ( w9534 , w9533 , w11004 );
not ( w9535 , w9534 );
and ( w9536 , w9535 , w8891 );
and ( w9537 , w9536 , w9551 );
nor ( w9538 , w9537 , w9133 );
and ( w9539 , w9439 , w9193 );
and ( w9540 , w9539 , w8891 );
and ( w9541 , w9540 , w10188 );
and ( w9542 , w9538 , w9554 );
not ( w9543 , w9542 );
and ( w9544 , w9543 , w8891 );
and ( w9545 , w9544 , w10188 );
nor ( w9546 , w9545 , w9027 );
nor ( w9547 , w9546 , w9241 );
nor ( w9548 , w9547 , w9012 );
not ( w9549 , w9548 );
and ( w9550 , w9549 , w8891 );
not ( w9551 , w9188 );
and ( w9552 , w9550 , w9551 );
nor ( w9553 , w9552 , w9133 );
not ( w9554 , w9541 );
and ( w9555 , w9553 , w9554 );
not ( w9556 , w9555 );
and ( w9557 , w9556 , w8891 );
and ( w9558 , w9557 , w10188 );
nor ( w9559 , w9558 , w9027 );
nor ( w9560 , w9020 , w9559 );
nor ( w9561 , w9560 , w9027 );
not ( w9562 , w9517 );
and ( w9563 , w9562 , w9561 );
and ( w9564 , w9563 , w9804 );
not ( w9565 , w9564 );
and ( w9566 , w9565 , w8891 );
and ( w9567 , w9566 , w10188 );
not ( w9568 , w9513 );
and ( w9569 , w9568 , w9567 );
and ( w9570 , w9569 , w8891 );
and ( w9571 , w9570 , w10188 );
and ( w9572 , w9571 , w8891 );
and ( w9573 , w10179 , w9572 );
nor ( w9574 , w9573 , w9285 );
and ( w9575 , w9574 , w9758 );
not ( w9576 , w9575 );
and ( w9577 , w9576 , w9567 );
nor ( w9578 , w9577 , w9027 );
and ( w9579 , w9490 , w9578 );
and ( w9580 , w9579 , w10615 );
and ( w9581 , w8895 , w9439 );
not ( w9582 , w9581 );
and ( w9583 , w9582 , w9578 );
and ( w9584 , w9583 , w9241 );
not ( w9585 , w9584 );
and ( w9586 , w9585 , w8891 );
nor ( w9587 , w9586 , w9285 );
and ( w9588 , w9587 , w9758 );
not ( w9589 , w9588 );
and ( w9590 , w9589 , w9567 );
and ( w9591 , w9590 , w8891 );
and ( w9592 , w9591 , w10188 );
nor ( w9593 , w9592 , w9027 );
nor ( w9594 , w9580 , w9593 );
and ( w9595 , w9594 , w8891 );
nor ( w9596 , w9595 , w9285 );
and ( w9597 , w9596 , w9758 );
not ( w9598 , w9597 );
and ( w9599 , w9598 , w9567 );
nor ( w9600 , w9599 , w9027 );
not ( w9601 , w8920 );
and ( w9602 , w9601 , w9600 );
nor ( w9603 , w9602 , w9593 );
and ( w9604 , w9603 , w8891 );
and ( w9605 , w9604 , w9567 );
not ( w9606 , w9605 );
and ( w9607 , w9480 , w9606 );
not ( w9608 , w9607 );
and ( w9609 , w9608 , w9567 );
nor ( w9610 , w9609 , w9027 );
nor ( w9611 , w9020 , w9610 );
nor ( w9612 , w9611 , w9285 );
and ( w9613 , w9612 , w9758 );
not ( w9614 , w9613 );
and ( w9615 , w9614 , w9567 );
nor ( w9616 , w9615 , w9027 );
not ( w9617 , w9474 );
and ( w9618 , w9617 , w9616 );
not ( w9619 , w9285 );
and ( w9620 , w9618 , w9619 );
and ( w9621 , w9620 , w9758 );
not ( w9622 , w9621 );
and ( w9623 , w9622 , w9567 );
nor ( w9624 , w9623 , w9027 );
not ( w9625 , w9463 );
and ( w9626 , w9625 , w9624 );
and ( w9627 , w9626 , w10905 );
nor ( w9628 , w9627 , w9020 );
not ( w9629 , w9628 );
and ( w9630 , w9629 , w8922 );
nor ( w9631 , w9630 , w9286 );
not ( w9632 , w9631 );
and ( w9633 , w9632 , w9624 );
and ( w9634 , w9633 , w8922 );
and ( w9635 , w9634 , w9624 );
and ( w9636 , w9635 , w8922 );
and ( w9637 , w9636 , w9935 );
and ( w9638 , w9637 , w8922 );
not ( w9639 , w9638 );
and ( w9640 , w9639 , w8891 );
not ( w9641 , w9640 );
and ( w9642 , w9641 , w8923 );
not ( w9643 , w9642 );
and ( w9644 , w9643 , w8879 );
and ( w9645 , w9644 , w8891 );
and ( w9646 , w8902 , w13206 );
and ( w9647 , w9439 , w10179 );
not ( w9648 , w9647 );
and ( w9649 , w9648 , w9633 );
and ( w9650 , w9649 , w8922 );
not ( w9651 , w9650 );
and ( w9652 , w9651 , w8909 );
nor ( w9653 , w9652 , w8905 );
and ( w9654 , w9653 , w8906 );
and ( w9655 , w9654 , w9241 );
not ( w9656 , w9655 );
and ( w9657 , w9656 , w8891 );
and ( w9658 , w9657 , w8890 );
and ( w9659 , w9658 , w8891 );
and ( w9660 , w9659 , w8893 );
not ( w9661 , w9660 );
and ( w9662 , w9661 , w9624 );
not ( w9663 , w9646 );
and ( w9664 , w9663 , w9662 );
not ( w9665 , w9664 );
and ( w9666 , w9665 , w8890 );
and ( w9667 , w9666 , w8891 );
and ( w9668 , w9667 , w8893 );
not ( w9669 , w9668 );
and ( w9670 , w9669 , w9624 );
and ( w9671 , w8890 , w9964 );
and ( w9672 , w9671 , w8891 );
and ( w9673 , w9672 , w8879 );
and ( w9674 , w9673 , w8891 );
and ( w9675 , w9636 , g39 );
and ( w9676 , w9675 , w8923 );
not ( w9677 , w9676 );
and ( w9678 , w9677 , w8879 );
not ( w9679 , w9678 );
and ( w9680 , w9679 , g13 );
and ( w9681 , w9680 , w9020 );
and ( w9682 , w9681 , w9028 );
and ( w9683 , w9682 , w8922 );
and ( w9684 , w9683 , w9624 );
and ( w9685 , w9684 , w10905 );
and ( w9686 , w9674 , w10008 );
and ( w9687 , w9686 , w8893 );
not ( w9688 , w9687 );
and ( w9689 , w9688 , w9624 );
not ( w9690 , w9689 );
and ( w9691 , w9645 , w9690 );
not ( w9692 , w9691 );
and ( w9693 , w9692 , w8922 );
and ( w9694 , w9693 , w9002 );
and ( w9695 , w8879 , g38 );
and ( w9696 , w9695 , g25 );
nor ( w9697 , w9696 , w9085 );
not ( w9698 , w9697 );
and ( w9699 , w9698 , w8891 );
and ( w9700 , w8879 , g44 );
and ( w9701 , w9700 , g27 );
nor ( w9702 , w9699 , w9701 );
not ( w9703 , w9702 );
and ( w9704 , w9703 , w8891 );
not ( w9705 , w9694 );
and ( w9706 , w9705 , w9704 );
not ( w9707 , w9706 );
and ( w9708 , w9707 , w9013 );
not ( w9709 , w9708 );
and ( w9710 , w9709 , w8891 );
nor ( w9711 , g38 , g25 );
and ( w9712 , w13511 , w8891 );
and ( w9713 , w9712 , w9085 );
nor ( w9714 , w9713 , w9696 );
not ( w9715 , w9714 );
and ( w9716 , w9715 , w8891 );
and ( w9717 , w9716 , w8879 );
and ( w9718 , w9717 , w9109 );
nor ( w9719 , w9718 , w9701 );
not ( w9720 , w9719 );
and ( w9721 , w9720 , w8879 );
and ( w9722 , w9721 , w8891 );
and ( w9723 , w9710 , w9722 );
and ( w9724 , w11760 , w8879 );
and ( w9725 , w9723 , w9724 );
and ( w9726 , w9725 , w9701 );
and ( w9727 , w8909 , w8891 );
not ( w9728 , w9727 );
and ( w9729 , w9728 , w8922 );
not ( w9730 , w9729 );
and ( w9731 , w9730 , w8879 );
and ( w9732 , w9731 , w10662 );
and ( w9733 , w9439 , w8909 );
not ( w9734 , w9733 );
and ( w9735 , w9734 , w8922 );
nor ( w9736 , w9085 , w9435 );
not ( w9737 , w9736 );
and ( w9738 , w9737 , w8891 );
nor ( w9739 , w9738 , w9704 );
not ( w9740 , w9739 );
and ( w9741 , w9740 , w8891 );
and ( w9742 , w9741 , w9113 );
not ( w9743 , w9742 );
and ( w9744 , w9743 , w8922 );
and ( w9745 , w8922 , g44 );
not ( w9746 , w9745 );
and ( w9747 , w9746 , w8879 );
not ( w9748 , w9747 );
and ( w9749 , w9748 , g27 );
not ( w9750 , w9749 );
and ( w9751 , w9750 , w9406 );
and ( w9752 , w9933 , w9002 );
nor ( w9753 , w9744 , w9752 );
and ( w9754 , w9753 , w8891 );
not ( w9755 , w9754 );
and ( w9756 , w9755 , w9013 );
and ( w9757 , w9735 , w9756 );
not ( w9758 , w9125 );
and ( w9759 , w9757 , w9758 );
and ( w9760 , w9759 , w9286 );
not ( w9761 , w8910 );
and ( w9762 , w9761 , w8879 );
and ( w9763 , w9762 , w8891 );
and ( w9764 , w8891 , w10949 );
nor ( w9765 , w9764 , w8909 );
not ( w9766 , w9765 );
and ( w9767 , w9766 , w9439 );
and ( w9768 , w9767 , w9435 );
and ( w9769 , w9768 , w8890 );
and ( w9770 , w9769 , w8891 );
nor ( w9771 , w9770 , w9085 );
not ( w9772 , w9696 );
and ( w9773 , w9771 , w9772 );
not ( w9774 , w9773 );
and ( w9775 , w9774 , w8891 );
and ( w9776 , w9775 , w8879 );
and ( w9777 , w9776 , w8891 );
nor ( w9778 , w9777 , w9701 );
not ( w9779 , w9778 );
and ( w9780 , w9779 , w8891 );
and ( w9781 , w9763 , w9780 );
and ( w9782 , w9781 , w8890 );
and ( w9783 , w9782 , w8879 );
and ( w9784 , w9783 , w8891 );
not ( w9785 , w9784 );
and ( w9786 , w9785 , w9627 );
nor ( w9787 , w9786 , w9286 );
and ( w9788 , w9787 , w8891 );
and ( w9789 , w9788 , w8890 );
and ( w9790 , w9789 , w8891 );
and ( w9791 , w9790 , w8893 );
not ( w9792 , w9791 );
and ( w9793 , w9792 , w9624 );
not ( w9794 , w9793 );
and ( w9795 , w8891 , w9794 );
and ( w9796 , w9795 , w8879 );
and ( w9797 , w9796 , w9113 );
not ( w9798 , w9797 );
and ( w9799 , w9798 , w8922 );
nor ( w9800 , w9799 , w9752 );
not ( w9801 , w9800 );
and ( w9802 , w9801 , w8922 );
and ( w9803 , w9802 , w9627 );
not ( w9804 , w9133 );
and ( w9805 , w9803 , w9804 );
not ( w9806 , w9805 );
and ( w9807 , w9806 , w8891 );
not ( w9808 , w9807 );
and ( w9809 , w9808 , w9013 );
and ( w9810 , w9809 , w8922 );
not ( w9811 , w9810 );
and ( w9812 , w9811 , w8891 );
nor ( w9813 , w9812 , w9249 );
not ( w9814 , w9813 );
and ( w9815 , w9814 , w8891 );
not ( w9816 , w9815 );
and ( w9817 , w9816 , w9028 );
and ( w9818 , w9817 , w8922 );
and ( w9819 , w9818 , w9624 );
nor ( w9820 , w9760 , w9819 );
and ( w9821 , w9820 , w10978 );
nor ( w9822 , w9821 , w9012 );
not ( w9823 , w9822 );
and ( w9824 , w9823 , w8891 );
and ( w9825 , w9824 , w8879 );
and ( w9826 , w9825 , w8891 );
and ( w9827 , w9826 , w11029 );
not ( w9828 , w9827 );
and ( w9829 , w9828 , w8922 );
and ( w9830 , w9829 , g36 );
not ( w9831 , w9830 );
and ( w9832 , w9831 , w8879 );
not ( w9833 , w9832 );
and ( w9834 , w9833 , g11 );
not ( w9835 , w9834 );
and ( w9836 , w9835 , w8891 );
not ( w9837 , w9836 );
and ( w9838 , w9837 , w9241 );
not ( w9839 , w9838 );
and ( w9840 , w9839 , w8891 );
and ( w9841 , w9439 , w8879 );
and ( w9842 , w9841 , g48 );
and ( w9843 , w9842 , g31 );
not ( w9844 , w9843 );
and ( w9845 , w9844 , w8922 );
and ( w9846 , w8922 , w10723 );
not ( w9847 , w9846 );
and ( w9848 , w9847 , w8891 );
and ( w9849 , w9848 , w8879 );
not ( w9850 , w9752 );
and ( w9851 , w9849 , w9850 );
not ( w9852 , w9851 );
and ( w9853 , w9852 , w9013 );
and ( w9854 , w9853 , w8923 );
and ( w9855 , w9854 , w9028 );
and ( w9856 , w9855 , w8922 );
not ( w9857 , w9856 );
and ( w9858 , w9857 , w8891 );
and ( w9859 , w9858 , w8893 );
not ( w9860 , w9859 );
and ( w9861 , w9860 , w9624 );
and ( w9862 , w9845 , w9861 );
nor ( w9863 , w9862 , w8997 );
and ( w9864 , w9863 , w8891 );
nor ( w9865 , w9864 , w9012 );
and ( w9866 , w9865 , w9478 );
not ( w9867 , w9866 );
and ( w9868 , w9867 , w9133 );
and ( w9869 , w9013 , w10723 );
not ( w9870 , w9869 );
and ( w9871 , w9870 , w8891 );
and ( w9872 , w9871 , w8879 );
not ( w9873 , w9872 );
and ( w9874 , w9873 , w8922 );
not ( w9875 , w9874 );
and ( w9876 , w9875 , w8891 );
and ( w9877 , w9751 , w10978 );
not ( w9878 , w9877 );
and ( w9879 , w9878 , w9002 );
and ( w9880 , w9879 , w9013 );
and ( w9881 , w9880 , w11004 );
not ( w9882 , w9881 );
and ( w9883 , w9882 , w8891 );
not ( w9884 , w9883 );
and ( w9885 , w9884 , w9028 );
and ( w9886 , w9885 , w8922 );
not ( w9887 , w9886 );
and ( w9888 , w9887 , w8891 );
and ( w9889 , w9888 , w8893 );
not ( w9890 , w9889 );
and ( w9891 , w9890 , w9624 );
and ( w9892 , w8922 , w9891 );
and ( w9893 , w9892 , w9627 );
nor ( w9894 , w9893 , w9286 );
not ( w9895 , w9894 );
and ( w9896 , w9895 , w8922 );
and ( w9897 , w9896 , w8923 );
not ( w9898 , w9897 );
and ( w9899 , w9898 , w8893 );
not ( w9900 , w9899 );
and ( w9901 , w9900 , w9624 );
not ( w9902 , w9901 );
and ( w9903 , w9876 , w9902 );
not ( w9904 , w9903 );
and ( w9905 , w9904 , w9627 );
nor ( w9906 , w9905 , w9286 );
not ( w9907 , w9906 );
and ( w9908 , w9907 , w8922 );
and ( w9909 , w9908 , w8923 );
and ( w9910 , w9909 , w9028 );
and ( w9911 , w9910 , w8922 );
not ( w9912 , w9911 );
and ( w9913 , w9912 , w8891 );
and ( w9914 , w9913 , w8893 );
not ( w9915 , w9914 );
and ( w9916 , w9915 , w9624 );
not ( w9917 , w9868 );
and ( w9918 , w9917 , w9916 );
and ( w9919 , w9918 , w8922 );
and ( w9920 , w9919 , w8923 );
not ( w9921 , w9920 );
and ( w9922 , w9921 , w8879 );
and ( w9923 , w9922 , w8891 );
nor ( w9924 , w9923 , w9193 );
not ( w9925 , w9924 );
and ( w9926 , w9925 , w8891 );
and ( w9927 , w9926 , w8893 );
not ( w9928 , w9927 );
and ( w9929 , w9928 , w9624 );
and ( w9930 , w9929 , w10905 );
and ( w9931 , w9840 , w9995 );
and ( w9932 , w9931 , w8891 );
not ( w9933 , w9751 );
and ( w9934 , w8922 , w9933 );
not ( w9935 , w9439 );
and ( w9936 , w9934 , w9935 );
not ( w9937 , w9936 );
and ( w9938 , w9937 , w8891 );
and ( w9939 , w9938 , w10978 );
not ( w9940 , w9939 );
and ( w9941 , w9940 , w9002 );
and ( w9942 , w9941 , w9013 );
not ( w9943 , w9942 );
and ( w9944 , w9943 , w8891 );
nor ( w9945 , w9944 , w9012 );
and ( w9946 , w9945 , w9478 );
not ( w9947 , w9946 );
and ( w9948 , w9947 , w9133 );
not ( w9949 , w9948 );
and ( w9950 , w9949 , w9901 );
and ( w9951 , w9950 , w8922 );
not ( w9952 , w9951 );
and ( w9953 , w9952 , w8891 );
and ( w9954 , w9953 , w8879 );
and ( w9955 , w9954 , w8891 );
not ( w9956 , w9955 );
and ( w9957 , w9956 , w8923 );
not ( w9958 , w9957 );
and ( w9959 , w9958 , w8879 );
and ( w9960 , w9959 , w8891 );
nor ( w9961 , w9960 , w9193 );
not ( w9962 , w9961 );
and ( w9963 , w9962 , w8891 );
not ( w9964 , w9670 );
and ( w9965 , w9963 , w9964 );
and ( w9966 , w9965 , w8891 );
not ( w9967 , w9966 );
and ( w9968 , w9967 , w9028 );
and ( w9969 , w9968 , w8922 );
not ( w9970 , w9969 );
and ( w9971 , w9970 , w8891 );
and ( w9972 , w9971 , w8893 );
not ( w9973 , w9972 );
and ( w9974 , w9973 , w9624 );
and ( w9975 , w9974 , w10905 );
not ( w9976 , w9975 );
and ( w9977 , w9932 , w9976 );
not ( w9978 , w9977 );
and ( w9979 , w9978 , w9028 );
and ( w9980 , w9979 , w8922 );
not ( w9981 , w9980 );
and ( w9982 , w9981 , w8893 );
not ( w9983 , w9982 );
and ( w9984 , w9983 , w9624 );
not ( w9985 , w9732 );
and ( w9986 , w9985 , w9984 );
and ( w9987 , w9986 , w8922 );
and ( w9988 , w9987 , g36 );
not ( w9989 , w9988 );
and ( w9990 , w9989 , w8879 );
not ( w9991 , w9990 );
and ( w9992 , w9991 , g11 );
not ( w9993 , w9992 );
and ( w9994 , w9993 , w8891 );
not ( w9995 , w9930 );
and ( w9996 , w9994 , w9995 );
and ( w9997 , w9996 , w8891 );
not ( w9998 , w9997 );
and ( w9999 , w9998 , w8922 );
not ( w10000 , w9999 );
and ( w10001 , w10000 , w8893 );
not ( w10002 , w10001 );
and ( w10003 , w10002 , w9624 );
not ( w10004 , w9726 );
and ( w10005 , w10004 , w10003 );
not ( w10006 , w10005 );
and ( w10007 , w10006 , w8891 );
not ( w10008 , w9685 );
and ( w10009 , w10007 , w10008 );
not ( w10010 , w10009 );
and ( w10011 , w10010 , w9028 );
and ( w10012 , w10011 , w8922 );
and ( w10013 , w10012 , w9624 );
and ( w10014 , w10013 , w10905 );
and ( w10015 , w9421 , w10138 );
nor ( w10016 , w9379 , w10015 );
and ( w10017 , w9406 , w10978 );
not ( w10018 , w9373 );
and ( w10019 , w8922 , w10018 );
and ( w10020 , w10052 , w10019 );
and ( w10021 , w10020 , w8865 );
and ( w10022 , w10021 , w8922 );
and ( w10023 , w10022 , w9002 );
nor ( w10024 , w10023 , w9008 );
not ( w10025 , w10024 );
and ( w10026 , w10025 , w9016 );
and ( w10027 , w10026 , w8865 );
and ( w10028 , w10027 , w13474 );
and ( w10029 , w10028 , w13477 );
not ( w10030 , w10029 );
and ( w10031 , w10030 , w8879 );
and ( w10032 , w10031 , w10138 );
not ( w10033 , w10016 );
and ( w10034 , w10033 , w10032 );
and ( w10035 , w10034 , w8879 );
not ( w10036 , w10035 );
and ( w10037 , w10036 , w8865 );
not ( w10038 , w10037 );
and ( w10039 , w10038 , g48 );
and ( w10040 , w10039 , g31 );
not ( w10041 , w10040 );
and ( w10042 , w10041 , w8922 );
not ( w10043 , w10015 );
and ( w10044 , w8923 , w10043 );
nor ( w10045 , w10044 , w10014 );
nor ( w10046 , w10045 , w9375 );
and ( w10047 , w10046 , g23 );
not ( w10048 , w10047 );
and ( w10049 , w10048 , w8891 );
and ( w10050 , w8923 , w10082 );
and ( w10051 , w8879 , w13204 );
not ( w10052 , w10017 );
and ( w10053 , w10052 , w8865 );
and ( w10054 , w10053 , w10019 );
and ( w10055 , w10054 , w8922 );
and ( w10056 , w10055 , w9002 );
nor ( w10057 , w10056 , w9008 );
and ( w10058 , w10057 , w13206 );
not ( w10059 , w10058 );
and ( w10060 , w10059 , w8865 );
and ( w10061 , w10060 , w13474 );
and ( w10062 , w10061 , w13477 );
not ( w10063 , w10062 );
and ( w10064 , w10063 , w8879 );
and ( w10065 , w10064 , w10138 );
and ( w10066 , w10051 , w10065 );
not ( w10067 , w10066 );
and ( w10068 , w10067 , w8865 );
and ( w10069 , w10068 , w9016 );
nor ( w10070 , w10069 , w10014 );
not ( w10071 , w10070 );
and ( w10072 , w8865 , w10071 );
and ( w10073 , w10072 , w10082 );
and ( w10074 , w10073 , w8865 );
and ( w10075 , w10074 , w13474 );
and ( w10076 , w10075 , w13477 );
not ( w10077 , w10076 );
and ( w10078 , w10077 , w8879 );
and ( w10079 , w10078 , w10138 );
not ( w10080 , w10079 );
and ( w10081 , w8922 , w10080 );
not ( w10082 , w10032 );
and ( w10083 , w10081 , w10082 );
and ( w10084 , w10083 , w8865 );
and ( w10085 , w10084 , w13474 );
and ( w10086 , w10085 , w13477 );
not ( w10087 , w10086 );
and ( w10088 , w10087 , w8879 );
and ( w10089 , w10088 , w10138 );
not ( w10090 , w10089 );
and ( w10091 , w8923 , w10090 );
nor ( w10092 , w10091 , w10014 );
not ( w10093 , w10050 );
and ( w10094 , w10093 , w10092 );
not ( w10095 , w10094 );
and ( w10096 , w10095 , w8922 );
and ( w10097 , w10096 , w8865 );
and ( w10098 , w10097 , w13474 );
and ( w10099 , w10098 , w13477 );
not ( w10100 , w10099 );
and ( w10101 , w10100 , w8879 );
and ( w10102 , w10101 , w10138 );
and ( w10103 , w10049 , w10102 );
not ( w10104 , w10103 );
and ( w10105 , w10104 , w8922 );
and ( w10106 , w10105 , w8865 );
and ( w10107 , w10106 , w13474 );
and ( w10108 , w10107 , w13477 );
not ( w10109 , w10108 );
and ( w10110 , w10109 , w8879 );
and ( w10111 , w10110 , w10138 );
and ( w10112 , w10042 , w10127 );
and ( w10113 , w10112 , w8865 );
and ( w10114 , w10113 , w13474 );
and ( w10115 , w10114 , w13477 );
not ( w10116 , w10115 );
and ( w10117 , w10116 , w8879 );
and ( w10118 , w10117 , w10138 );
not ( w10119 , w10118 );
and ( w10120 , w8923 , w10119 );
not ( w10121 , w10120 );
and ( w10122 , w10121 , w8879 );
and ( w10123 , w10122 , g48 );
and ( w10124 , w10123 , g31 );
not ( w10125 , w10124 );
and ( w10126 , w10125 , w8922 );
not ( w10127 , w10111 );
and ( w10128 , w10126 , w10127 );
nor ( w10129 , w10128 , w10014 );
not ( w10130 , w9021 );
and ( w10131 , w10130 , w10129 );
not ( w10132 , w10131 );
and ( w10133 , w10132 , w8865 );
and ( w10134 , w10133 , w13474 );
and ( w10135 , w10134 , w13477 );
not ( w10136 , w10135 );
and ( w10137 , w10136 , w8879 );
not ( w10138 , w10014 );
and ( w10139 , w10137 , w10138 );
and ( w10140 , w9360 , w10139 );
not ( w10141 , w9350 );
and ( w10142 , w10141 , w10140 );
and ( w10143 , w10142 , w8891 );
and ( w10144 , w10143 , w10188 );
and ( w10145 , w10144 , w10234 );
and ( w10146 , w10145 , w8891 );
and ( w10147 , w10146 , w10139 );
not ( w10148 , w9325 );
and ( w10149 , w10148 , w10147 );
and ( w10150 , w10149 , w9303 );
and ( w10151 , w10150 , w10200 );
nor ( w10152 , w8920 , w9520 );
nor ( w10153 , w10152 , w9525 );
and ( w10154 , w10153 , w10179 );
nor ( w10155 , w10154 , w9193 );
not ( w10156 , w10155 );
and ( w10157 , w10156 , w9122 );
and ( w10158 , w10157 , w9244 );
and ( w10159 , w10158 , w8891 );
and ( w10160 , w10159 , w10179 );
not ( w10161 , w10160 );
and ( w10162 , w10161 , w8922 );
and ( w10163 , w10162 , w8865 );
nor ( w10164 , w10163 , w9286 );
nor ( w10165 , w10151 , w10164 );
and ( w10166 , w10165 , w11004 );
not ( w10167 , w10166 );
and ( w10168 , w10167 , w8891 );
and ( w10169 , w10168 , w9122 );
nor ( w10170 , w10169 , w8988 );
nor ( w10171 , w10170 , w9188 );
not ( w10172 , w10171 );
and ( w10173 , w10172 , w8922 );
and ( w10174 , w10173 , w8923 );
and ( w10175 , w10174 , w10615 );
not ( w10176 , w10175 );
and ( w10177 , w10176 , w9244 );
and ( w10178 , w10177 , w8891 );
not ( w10179 , w9020 );
and ( w10180 , w10178 , w10179 );
not ( w10181 , w10180 );
and ( w10182 , w10181 , w8922 );
and ( w10183 , w10182 , w8865 );
and ( w10184 , w10183 , w8933 );
not ( w10185 , w10184 );
and ( w10186 , w10185 , w10140 );
and ( w10187 , w10186 , w8891 );
not ( w10188 , w9237 );
and ( w10189 , w10187 , w10188 );
and ( w10190 , w10189 , w10234 );
and ( w10191 , w10190 , w8891 );
and ( w10192 , w10191 , w10139 );
nor ( w10193 , w9322 , w10192 );
and ( w10194 , w10193 , w8933 );
not ( w10195 , w10194 );
and ( w10196 , w10195 , w10140 );
and ( w10197 , w10196 , w10234 );
not ( w10198 , w9158 );
and ( w10199 , w10198 , w10197 );
not ( w10200 , w9205 );
and ( w10201 , w10199 , w10200 );
not ( w10202 , w10201 );
and ( w10203 , w10202 , w8865 );
and ( w10204 , w10203 , w10994 );
not ( w10205 , w10204 );
and ( w10206 , w10205 , w8879 );
and ( w10207 , w10206 , w8891 );
and ( w10208 , w10207 , w10999 );
not ( w10209 , w10208 );
and ( w10210 , w10209 , w8865 );
and ( w10211 , w10210 , w10276 );
nor ( w10212 , w10211 , w8997 );
not ( w10213 , w10212 );
and ( w10214 , w10213 , w8865 );
and ( w10215 , w10214 , w8922 );
and ( w10216 , w10215 , w9002 );
nor ( w10217 , w10216 , w9008 );
not ( w10218 , w10217 );
and ( w10219 , w10218 , w8922 );
and ( w10220 , w10219 , w8923 );
and ( w10221 , w10220 , w9016 );
nor ( w10222 , w10221 , w9021 );
not ( w10223 , w10222 );
and ( w10224 , w10223 , w8865 );
and ( w10225 , w10224 , w8922 );
nor ( w10226 , w10225 , w9241 );
nor ( w10227 , w10226 , w9122 );
not ( w10228 , w10227 );
and ( w10229 , w10228 , w9027 );
nor ( w10230 , w10229 , w10192 );
and ( w10231 , w10230 , w8933 );
not ( w10232 , w10231 );
and ( w10233 , w10232 , w10140 );
not ( w10234 , w9286 );
and ( w10235 , w10233 , w10234 );
and ( w10236 , w10235 , w8891 );
and ( w10237 , w10236 , w10139 );
not ( w10238 , w10237 );
and ( w10239 , w8865 , w10238 );
and ( w10240 , w10239 , w10994 );
not ( w10241 , w10240 );
and ( w10242 , w10241 , w8879 );
and ( w10243 , w10242 , w8891 );
and ( w10244 , w10243 , w10999 );
not ( w10245 , w10244 );
and ( w10246 , w10245 , w8865 );
and ( w10247 , w10246 , w10276 );
nor ( w10248 , w10247 , w8997 );
not ( w10249 , w10248 );
and ( w10250 , w10249 , w8865 );
and ( w10251 , w10250 , w8922 );
and ( w10252 , w10251 , w9002 );
nor ( w10253 , w10252 , w9008 );
not ( w10254 , w10253 );
and ( w10255 , w10254 , w8922 );
and ( w10256 , w10255 , w8923 );
and ( w10257 , w10256 , w9016 );
nor ( w10258 , w10257 , w9021 );
not ( w10259 , w10258 );
and ( w10260 , w10259 , w8865 );
and ( w10261 , w10260 , w8922 );
nor ( w10262 , w10261 , w9241 );
nor ( w10263 , w10262 , w9122 );
not ( w10264 , w10263 );
and ( w10265 , w10264 , w9027 );
nor ( w10266 , w10265 , w10192 );
nor ( w10267 , w10266 , w9286 );
nor ( w10268 , w9157 , w10267 );
and ( w10269 , w8906 , w10268 );
and ( w10270 , w10269 , w10329 );
not ( w10271 , w10270 );
and ( w10272 , w10271 , w8890 );
and ( w10273 , w10272 , w8891 );
and ( w10274 , w10273 , w8879 );
and ( w10275 , w10274 , w10662 );
not ( w10276 , w8994 );
and ( w10277 , w8922 , w10276 );
not ( w10278 , w10277 );
and ( w10279 , w10278 , w8879 );
and ( w10280 , w10279 , w8891 );
not ( w10281 , w10280 );
and ( w10282 , w10281 , w9013 );
and ( w10283 , w10282 , w11004 );
and ( w10284 , w10283 , w9002 );
and ( w10285 , w10284 , w10568 );
not ( w10286 , w10285 );
and ( w10287 , w10286 , w8891 );
nor ( w10288 , w10287 , w9193 );
not ( w10289 , w10288 );
and ( w10290 , w10289 , w8891 );
and ( w10291 , w10290 , w8879 );
and ( w10292 , w10291 , w8891 );
and ( w10293 , w8891 , w8936 );
nor ( w10294 , w10293 , w8994 );
not ( w10295 , w10294 );
and ( w10296 , w10295 , w8891 );
and ( w10297 , w10296 , w10949 );
not ( w10298 , w10297 );
and ( w10299 , w10298 , w10268 );
and ( w10300 , w10299 , w10329 );
nor ( w10301 , w8936 , w9224 );
nor ( w10302 , w10300 , w10301 );
and ( w10303 , w10302 , w8891 );
nor ( w10304 , w10303 , w8988 );
and ( w10305 , w9153 , w8906 );
and ( w10306 , w10393 , w8890 );
nor ( w10307 , w10306 , w8909 );
not ( w10308 , w10307 );
and ( w10309 , w10308 , w8879 );
and ( w10310 , w10309 , w8891 );
and ( w10311 , w10310 , w8890 );
not ( w10312 , w10311 );
and ( w10313 , w10312 , w8922 );
not ( w10314 , w10313 );
and ( w10315 , w10314 , w8891 );
and ( w10316 , w10315 , w8893 );
nor ( w10317 , w10316 , w10267 );
nor ( w10318 , w10304 , w10317 );
and ( w10319 , w10318 , w8890 );
and ( w10320 , w10319 , w8891 );
and ( w10321 , w10320 , w8893 );
nor ( w10322 , w10321 , w10267 );
not ( w10323 , w10322 );
and ( w10324 , w10323 , w8891 );
nor ( w10325 , w10324 , w9012 );
not ( w10326 , w10325 );
and ( w10327 , w10326 , w8879 );
and ( w10328 , w10327 , w8891 );
not ( w10329 , w8909 );
and ( w10330 , w10305 , w10329 );
not ( w10331 , w10330 );
and ( w10332 , w10331 , w8891 );
and ( w10333 , w10332 , w8890 );
not ( w10334 , w10333 );
and ( w10335 , w10334 , w8922 );
not ( w10336 , w10335 );
and ( w10337 , w10336 , w8891 );
and ( w10338 , w10337 , w8893 );
nor ( w10339 , w10338 , w10267 );
not ( w10340 , w10339 );
and ( w10341 , w10328 , w10340 );
not ( w10342 , w10317 );
and ( w10343 , w10341 , w10342 );
and ( w10344 , w10343 , w8891 );
and ( w10345 , w10344 , w8879 );
and ( w10346 , w10345 , w8891 );
nor ( w10347 , w9012 , w9224 );
not ( w10348 , w10347 );
and ( w10349 , w10348 , w8891 );
and ( w10350 , w10346 , w10349 );
and ( w10351 , w10350 , w8891 );
and ( w10352 , w9002 , w8865 );
not ( w10353 , w10352 );
and ( w10354 , w10353 , w8891 );
and ( w10355 , w10354 , w8879 );
and ( w10356 , w10355 , w9113 );
not ( w10357 , w10356 );
and ( w10358 , w10357 , w8922 );
and ( w10359 , w10358 , w8923 );
nor ( w10360 , w10359 , w9458 );
not ( w10361 , w10360 );
and ( w10362 , w8922 , w10361 );
and ( w10363 , w10362 , w9002 );
and ( w10364 , w10363 , w8922 );
nor ( w10365 , w10364 , w9241 );
and ( w10366 , w8922 , w10805 );
and ( w10367 , w10366 , w9002 );
nor ( w10368 , w10367 , w10317 );
not ( w10369 , w10368 );
and ( w10370 , w10369 , w8922 );
not ( w10371 , w10370 );
and ( w10372 , w10371 , w8891 );
and ( w10373 , w10372 , w9193 );
nor ( w10374 , w10373 , w9027 );
not ( w10375 , w10374 );
and ( w10376 , w10375 , w9122 );
and ( w10377 , w10376 , w8891 );
and ( w10378 , w10377 , w8879 );
and ( w10379 , w10378 , w8891 );
and ( w10380 , w10379 , w11029 );
not ( w10381 , w10380 );
and ( w10382 , w10381 , w8922 );
and ( w10383 , w10382 , w9039 );
and ( w10384 , w10383 , w8922 );
and ( w10385 , w10384 , w8928 );
and ( w10386 , w10385 , w8922 );
and ( w10387 , w10386 , w8865 );
and ( w10388 , w10387 , w8933 );
and ( w10389 , w10388 , w10994 );
not ( w10390 , w10389 );
and ( w10391 , w10390 , w8879 );
and ( w10392 , w10391 , w8891 );
not ( w10393 , w10305 );
and ( w10394 , w10393 , w8891 );
nor ( w10395 , w10394 , w8909 );
not ( w10396 , w10395 );
and ( w10397 , w10396 , w8891 );
and ( w10398 , w8890 , w10397 );
and ( w10399 , w10398 , w8879 );
and ( w10400 , w10399 , w8891 );
and ( w10401 , w10397 , w10139 );
and ( w10402 , w10401 , w8890 );
not ( w10403 , w10402 );
and ( w10404 , w10403 , w8922 );
not ( w10405 , w10404 );
and ( w10406 , w10405 , w8891 );
and ( w10407 , w10406 , w8893 );
nor ( w10408 , w10407 , w10267 );
not ( w10409 , w10408 );
and ( w10410 , w10409 , w8891 );
and ( w10411 , w10410 , w10139 );
and ( w10412 , w10400 , w10411 );
and ( w10413 , w10412 , w8985 );
not ( w10414 , w8977 );
and ( w10415 , w10414 , w8922 );
not ( w10416 , w10415 );
and ( w10417 , w10416 , w10397 );
and ( w10418 , w10417 , w8891 );
not ( w10419 , w10418 );
and ( w10420 , w10419 , w8928 );
and ( w10421 , w10420 , w8922 );
and ( w10422 , w10421 , w8933 );
not ( w10423 , w10422 );
and ( w10424 , w10423 , w10401 );
and ( w10425 , w10424 , w9214 );
not ( w10426 , w10425 );
and ( w10427 , w10426 , w8922 );
and ( w10428 , w8922 , w12962 );
and ( w10429 , w10428 , w12964 );
not ( w10430 , w10429 );
and ( w10431 , w10430 , w8879 );
not ( w10432 , w10427 );
and ( w10433 , w10432 , w10431 );
not ( w10434 , w10433 );
and ( w10435 , w10434 , w8922 );
not ( w10436 , w10435 );
and ( w10437 , w10436 , w8985 );
not ( w10438 , w10437 );
and ( w10439 , w10438 , w8865 );
and ( w10440 , w10439 , w8922 );
not ( w10441 , w10440 );
and ( w10442 , w10441 , w8891 );
not ( w10443 , w10442 );
and ( w10444 , w10443 , w9013 );
and ( w10445 , w10444 , w8865 );
not ( w10446 , w10445 );
and ( w10447 , w10446 , w9085 );
and ( w10448 , w10447 , w9724 );
nor ( w10449 , w9749 , w8989 );
not ( w10450 , w10449 );
and ( w10451 , w10450 , w8865 );
nor ( w10452 , w9696 , w9701 );
nor ( w10453 , w10451 , w10452 );
not ( w10454 , w10453 );
and ( w10455 , w10454 , w8922 );
and ( w10456 , w10455 , w9002 );
not ( w10457 , w10456 );
and ( w10458 , w10457 , w8891 );
and ( w10459 , w10458 , w9109 );
not ( w10460 , w10459 );
and ( w10461 , w10460 , w8922 );
and ( w10462 , w10461 , w9013 );
not ( w10463 , w10462 );
and ( w10464 , w10463 , w9724 );
not ( w10465 , w10464 );
and ( w10466 , w10465 , w8922 );
not ( w10467 , w10448 );
and ( w10468 , w10467 , w10466 );
and ( w10469 , w10468 , w9002 );
not ( w10470 , w10469 );
and ( w10471 , w10470 , w8891 );
and ( w10472 , w10471 , w10978 );
and ( w10473 , w10472 , w8890 );
not ( w10474 , w10473 );
and ( w10475 , w10474 , w8922 );
not ( w10476 , w10475 );
and ( w10477 , w10476 , w8891 );
and ( w10478 , w10477 , w8893 );
nor ( w10479 , w10478 , w10267 );
not ( w10480 , w10479 );
and ( w10481 , w10480 , w8891 );
and ( w10482 , w10481 , w10139 );
and ( w10483 , w9085 , w10482 );
not ( w10484 , w10483 );
and ( w10485 , w10484 , w10466 );
nor ( w10486 , w10485 , w10317 );
not ( w10487 , w10486 );
and ( w10488 , w10487 , w8922 );
and ( w10489 , w10488 , w10805 );
not ( w10490 , w10413 );
and ( w10491 , w10490 , w10489 );
not ( w10492 , w10491 );
and ( w10493 , w10492 , w8891 );
and ( w10494 , w10493 , w10978 );
not ( w10495 , w10494 );
and ( w10496 , w10495 , w8922 );
not ( w10497 , w10496 );
and ( w10498 , w10497 , w8890 );
not ( w10499 , w10498 );
and ( w10500 , w10499 , w8922 );
not ( w10501 , w10500 );
and ( w10502 , w10501 , w8891 );
and ( w10503 , w10502 , w8893 );
nor ( w10504 , w10503 , w10267 );
not ( w10505 , w10504 );
and ( w10506 , w10505 , w8891 );
and ( w10507 , w10506 , w10139 );
not ( w10508 , w9059 );
and ( w10509 , w10507 , w10508 );
not ( w10510 , w8970 );
and ( w10511 , w10509 , w10510 );
and ( w10512 , w10511 , w10969 );
not ( w10513 , w10512 );
and ( w10514 , w10513 , w8922 );
and ( w10515 , w10514 , w10322 );
and ( w10516 , w10515 , w10987 );
not ( w10517 , w10516 );
and ( w10518 , w10517 , w8891 );
not ( w10519 , w10518 );
and ( w10520 , w10519 , w8865 );
and ( w10521 , w10520 , w8933 );
not ( w10522 , w10521 );
and ( w10523 , w10522 , w10401 );
and ( w10524 , w10523 , w8985 );
nor ( w10525 , w10482 , w8988 );
nor ( w10526 , w10525 , w9059 );
and ( w10527 , w10526 , w10969 );
not ( w10528 , w10527 );
and ( w10529 , w10528 , w8928 );
and ( w10530 , w10529 , w8922 );
and ( w10531 , w10530 , w8933 );
not ( w10532 , w10531 );
and ( w10533 , w10532 , w10401 );
and ( w10534 , w10533 , w10999 );
not ( w10535 , w10534 );
and ( w10536 , w10535 , w8922 );
not ( w10537 , w10536 );
and ( w10538 , w10537 , w8985 );
not ( w10539 , w10538 );
and ( w10540 , w10539 , w8865 );
and ( w10541 , w10540 , w8922 );
and ( w10542 , w10541 , w8865 );
and ( w10543 , w10542 , w10466 );
not ( w10544 , w10543 );
and ( w10545 , w10544 , w8891 );
and ( w10546 , w10545 , w10978 );
not ( w10547 , w10546 );
and ( w10548 , w10547 , w10366 );
and ( w10549 , w10548 , w9002 );
nor ( w10550 , w10549 , w10317 );
and ( w10551 , w10550 , w8890 );
not ( w10552 , w10551 );
and ( w10553 , w10552 , w8922 );
not ( w10554 , w10553 );
and ( w10555 , w10554 , w8891 );
and ( w10556 , w10555 , w8893 );
nor ( w10557 , w10556 , w10267 );
not ( w10558 , w10557 );
and ( w10559 , w10558 , w8891 );
and ( w10560 , w10559 , w10139 );
nor ( w10561 , w10524 , w10560 );
not ( w10562 , w10561 );
and ( w10563 , w10562 , w8891 );
and ( w10564 , w10563 , w10978 );
not ( w10565 , w10564 );
and ( w10566 , w10565 , w10366 );
and ( w10567 , w10566 , w9002 );
not ( w10568 , w8988 );
and ( w10569 , w10567 , w10568 );
nor ( w10570 , w10569 , w10317 );
not ( w10571 , w10570 );
and ( w10572 , w10571 , w9013 );
and ( w10573 , w10572 , w11004 );
nor ( w10574 , w10573 , w10339 );
and ( w10575 , w10574 , w8891 );
and ( w10576 , w9846 , w9013 );
not ( w10577 , w10576 );
and ( w10578 , w10577 , w8891 );
and ( w10579 , w10578 , w8879 );
not ( w10580 , w10579 );
and ( w10581 , w10580 , w8923 );
nor ( w10582 , w10581 , w9458 );
not ( w10583 , w10582 );
and ( w10584 , w10583 , w8922 );
not ( w10585 , w10584 );
and ( w10586 , w10575 , w10585 );
and ( w10587 , w10586 , w8891 );
and ( w10588 , w10587 , w8879 );
and ( w10589 , w10588 , w8891 );
not ( w10590 , w10589 );
and ( w10591 , w10590 , w9241 );
not ( w10592 , w10591 );
and ( w10593 , w10592 , w8891 );
and ( w10594 , w10593 , w11029 );
and ( w10595 , w8989 , w8865 );
nor ( w10596 , w10595 , w8997 );
not ( w10597 , w10596 );
and ( w10598 , w10597 , w8922 );
and ( w10599 , w10598 , w8865 );
and ( w10600 , w10599 , w8922 );
and ( w10601 , w10600 , w9002 );
not ( w10602 , w10601 );
and ( w10603 , w10602 , w8891 );
and ( w10604 , w10603 , w8879 );
and ( w10605 , w10604 , w9113 );
not ( w10606 , w10605 );
and ( w10607 , w10606 , w8922 );
and ( w10608 , w10607 , w9013 );
and ( w10609 , w10608 , w8922 );
not ( w10610 , w10609 );
and ( w10611 , w10610 , w8891 );
and ( w10612 , w9186 , w8879 );
and ( w10613 , w10612 , w9113 );
nor ( w10614 , w10611 , w10613 );
not ( w10615 , w9193 );
and ( w10616 , w10614 , w10615 );
and ( w10617 , w10616 , w8922 );
not ( w10618 , w10617 );
and ( w10619 , w10618 , w9122 );
not ( w10620 , w10619 );
and ( w10621 , w10620 , w8922 );
and ( w10622 , w10621 , w8865 );
and ( w10623 , w10622 , w11022 );
and ( w10624 , w10623 , w8922 );
not ( w10625 , w10624 );
and ( w10626 , w10625 , w8891 );
and ( w10627 , w10626 , w8893 );
nor ( w10628 , w10627 , w10267 );
nor ( w10629 , w10628 , w9286 );
and ( w10630 , w10594 , w10629 );
not ( w10631 , w10630 );
and ( w10632 , w10631 , w8922 );
and ( w10633 , w10632 , w8865 );
not ( w10634 , w10633 );
and ( w10635 , w10634 , w8891 );
nor ( w10636 , w10635 , w9249 );
not ( w10637 , w10636 );
and ( w10638 , w10637 , w8891 );
and ( w10639 , w10638 , w8890 );
not ( w10640 , w10639 );
and ( w10641 , w10640 , w8922 );
not ( w10642 , w10641 );
and ( w10643 , w10642 , w8891 );
and ( w10644 , w10643 , w8893 );
nor ( w10645 , w10644 , w10267 );
not ( w10646 , w10645 );
and ( w10647 , w10646 , w8891 );
and ( w10648 , w10647 , w10139 );
nor ( w10649 , w10275 , w10648 );
not ( w10650 , w10649 );
and ( w10651 , w10650 , w9122 );
not ( w10652 , w10651 );
and ( w10653 , w10652 , w8922 );
and ( w10654 , w10653 , w8865 );
not ( w10655 , w10654 );
and ( w10656 , w10655 , w8891 );
and ( w10657 , w10656 , w8890 );
and ( w10658 , w10657 , w8891 );
and ( w10659 , w10658 , w8893 );
nor ( w10660 , w10659 , w10267 );
nor ( w10661 , w10660 , w9286 );
not ( w10662 , w8923 );
and ( w10663 , w10661 , w10662 );
nor ( w10664 , w10663 , w9027 );
and ( w10665 , w11039 , w10648 );
nor ( w10666 , w10665 , w9027 );
not ( w10667 , w10666 );
and ( w10668 , w10667 , w9122 );
not ( w10669 , w10668 );
and ( w10670 , w10669 , w8922 );
and ( w10671 , w10670 , w10805 );
not ( w10672 , w10671 );
and ( w10673 , w10672 , w8891 );
and ( w10674 , w10673 , w10139 );
not ( w10675 , w10674 );
and ( w10676 , w10664 , w10675 );
not ( w10677 , w10676 );
and ( w10678 , w10677 , w9122 );
and ( w10679 , w8865 , w9021 );
not ( w10680 , w9178 );
and ( w10681 , w10680 , w8922 );
and ( w10682 , w10681 , w8865 );
and ( w10683 , w10682 , w8923 );
and ( w10684 , w10683 , w9016 );
and ( w10685 , w10684 , w8922 );
nor ( w10686 , w10685 , w9241 );
nor ( w10687 , w10686 , w9122 );
not ( w10688 , w10687 );
and ( w10689 , w10688 , w9027 );
not ( w10690 , w10689 );
and ( w10691 , w10690 , w8865 );
and ( w10692 , w10691 , w11022 );
nor ( w10693 , w10679 , w10692 );
not ( w10694 , w10693 );
and ( w10695 , w10694 , w8865 );
and ( w10696 , w10695 , w8922 );
not ( w10697 , w10678 );
and ( w10698 , w10697 , w10696 );
and ( w10699 , w10698 , w8865 );
not ( w10700 , w10699 );
and ( w10701 , w10700 , w8891 );
and ( w10702 , w10701 , w8893 );
nor ( w10703 , w10702 , w10267 );
nor ( w10704 , w10703 , w9286 );
and ( w10705 , w10704 , w8891 );
and ( w10706 , w10705 , w10139 );
and ( w10707 , w10392 , w10706 );
not ( w10708 , w10707 );
and ( w10709 , w10708 , w8922 );
and ( w10710 , w10709 , w10805 );
not ( w10711 , w10710 );
and ( w10712 , w10711 , w8891 );
and ( w10713 , w10712 , w10139 );
nor ( w10714 , w10365 , w10713 );
and ( w10715 , w10714 , w9013 );
not ( w10716 , w10715 );
and ( w10717 , w10716 , w9724 );
and ( w10718 , w10717 , w8891 );
and ( w10719 , w10718 , w8879 );
and ( w10720 , w10719 , w8891 );
and ( w10721 , w10584 , w9013 );
and ( w10722 , w10721 , w11004 );
not ( w10723 , w9113 );
and ( w10724 , w10722 , w10723 );
not ( w10725 , w10724 );
and ( w10726 , w10725 , w8891 );
nor ( w10727 , w10726 , w9249 );
not ( w10728 , w10727 );
and ( w10729 , w10728 , w8891 );
and ( w10730 , w10729 , w8879 );
and ( w10731 , w10730 , w8891 );
and ( w10732 , w10731 , w11029 );
not ( w10733 , w10732 );
and ( w10734 , w10733 , w8922 );
and ( w10735 , w10734 , w10805 );
and ( w10736 , w10720 , w10797 );
nor ( w10737 , w10736 , w9249 );
not ( w10738 , w10737 );
and ( w10739 , w10738 , w8891 );
nor ( w10740 , w10739 , w9027 );
not ( w10741 , w10740 );
and ( w10742 , w10741 , w9122 );
and ( w10743 , w10742 , w8891 );
and ( w10744 , w10743 , w8879 );
and ( w10745 , w10744 , w8891 );
and ( w10746 , w10745 , w11029 );
not ( w10747 , w10746 );
and ( w10748 , w10747 , w8922 );
and ( w10749 , w10748 , w9039 );
and ( w10750 , w10749 , w8922 );
and ( w10751 , w10750 , w8928 );
and ( w10752 , w10751 , w8922 );
and ( w10753 , w10752 , w8865 );
and ( w10754 , w10753 , w8933 );
and ( w10755 , w10754 , w10994 );
not ( w10756 , w10755 );
and ( w10757 , w10756 , w8879 );
and ( w10758 , w10757 , w8891 );
and ( w10759 , w10758 , w10706 );
not ( w10760 , w10759 );
and ( w10761 , w10760 , w8922 );
and ( w10762 , w10761 , w10805 );
nor ( w10763 , w10762 , w9286 );
and ( w10764 , w10763 , w8891 );
and ( w10765 , w10764 , w10139 );
nor ( w10766 , w10351 , w10765 );
nor ( w10767 , w10766 , w10735 );
and ( w10768 , w10767 , w8891 );
nor ( w10769 , w10768 , w9027 );
not ( w10770 , w10769 );
and ( w10771 , w10770 , w9122 );
and ( w10772 , w10771 , w8891 );
and ( w10773 , w10772 , w8879 );
and ( w10774 , w10773 , w8891 );
and ( w10775 , w10774 , w11029 );
not ( w10776 , w10775 );
and ( w10777 , w10776 , w8922 );
and ( w10778 , w10852 , w8865 );
and ( w10779 , w10777 , w10778 );
and ( w10780 , w10779 , w10987 );
not ( w10781 , w10780 );
and ( w10782 , w10781 , w8891 );
not ( w10783 , w10782 );
and ( w10784 , w10783 , w8865 );
and ( w10785 , w10784 , w8933 );
and ( w10786 , w10785 , w10994 );
not ( w10787 , w10786 );
and ( w10788 , w10787 , w8879 );
and ( w10789 , w10788 , w8891 );
and ( w10790 , w10789 , w10706 );
and ( w10791 , w10790 , w8893 );
nor ( w10792 , w10791 , w10267 );
not ( w10793 , w10792 );
and ( w10794 , w10793 , w8891 );
and ( w10795 , w10794 , w10139 );
and ( w10796 , w10292 , w10795 );
not ( w10797 , w10735 );
and ( w10798 , w10796 , w10797 );
nor ( w10799 , w10798 , w9249 );
and ( w10800 , w9035 , w10905 );
not ( w10801 , w10800 );
and ( w10802 , w10801 , w9122 );
not ( w10803 , w10802 );
and ( w10804 , w10803 , w8922 );
not ( w10805 , w10267 );
and ( w10806 , w10804 , w10805 );
nor ( w10807 , w10799 , w10806 );
nor ( w10808 , w10807 , w9027 );
not ( w10809 , w10808 );
and ( w10810 , w10809 , w8891 );
and ( w10811 , w10810 , w9122 );
and ( w10812 , w10811 , w8891 );
and ( w10813 , w10812 , w8879 );
and ( w10814 , w10813 , w8891 );
and ( w10815 , w10814 , w11029 );
not ( w10816 , w10815 );
and ( w10817 , w10816 , w8922 );
and ( w10818 , w10817 , w10778 );
and ( w10819 , w10818 , w9039 );
and ( w10820 , w10819 , w10987 );
and ( w10821 , w10820 , w8922 );
not ( w10822 , w10821 );
and ( w10823 , w10822 , w8891 );
not ( w10824 , w10823 );
and ( w10825 , w10824 , w8928 );
and ( w10826 , w10825 , w8922 );
and ( w10827 , w10826 , w8865 );
and ( w10828 , w10827 , w8933 );
and ( w10829 , w10828 , w10994 );
not ( w10830 , w10829 );
and ( w10831 , w10830 , w8879 );
and ( w10832 , w10831 , w8891 );
and ( w10833 , w10832 , w10706 );
not ( w10834 , w10833 );
and ( w10835 , w10834 , w8922 );
not ( w10836 , w10835 );
and ( w10837 , w10836 , w8891 );
and ( w10838 , w10837 , w8893 );
nor ( w10839 , w10838 , w10267 );
nor ( w10840 , w10839 , w9286 );
and ( w10841 , w10840 , w8891 );
and ( w10842 , w10841 , w10139 );
nor ( w10843 , w10275 , w10842 );
not ( w10844 , w10843 );
and ( w10845 , w10844 , w9122 );
and ( w10846 , w10845 , w8890 );
and ( w10847 , w10846 , w8891 );
and ( w10848 , w10847 , w8893 );
nor ( w10849 , w10848 , w10267 );
nor ( w10850 , w10849 , w9286 );
nor ( w10851 , w9151 , w10850 );
not ( w10852 , w8978 );
and ( w10853 , w10851 , w10852 );
and ( w10854 , w10853 , w8922 );
and ( w10855 , w10854 , w8928 );
and ( w10856 , w10855 , w8865 );
and ( w10857 , w10856 , w8933 );
and ( w10858 , w10857 , w10994 );
not ( w10859 , w10858 );
and ( w10860 , w10859 , w8879 );
and ( w10861 , w10860 , w8891 );
and ( w10862 , w10861 , w10706 );
not ( w10863 , w10862 );
and ( w10864 , w10863 , w8865 );
not ( w10865 , w10864 );
and ( w10866 , w10865 , w8891 );
and ( w10867 , w10866 , w8893 );
nor ( w10868 , w10867 , w10267 );
nor ( w10869 , w10868 , w9286 );
and ( w10870 , w10869 , w8891 );
and ( w10871 , w10870 , w10139 );
nor ( w10872 , w9135 , w10871 );
not ( w10873 , w10872 );
and ( w10874 , w10873 , w8891 );
and ( w10875 , w10874 , w10139 );
not ( w10876 , w10875 );
and ( w10877 , w8922 , w10876 );
and ( w10878 , w10877 , w11046 );
not ( w10879 , w10878 );
and ( w10880 , w10879 , w8890 );
not ( w10881 , w10880 );
and ( w10882 , w10881 , w8922 );
not ( w10883 , w10882 );
and ( w10884 , w10883 , w8891 );
and ( w10885 , w10884 , w8893 );
nor ( w10886 , w9265 , w8989 );
and ( w10887 , w10886 , w10978 );
nor ( w10888 , w10887 , w8988 );
nor ( w10889 , w10888 , w9241 );
and ( w10890 , w10889 , w8891 );
and ( w10891 , w10890 , w8879 );
and ( w10892 , w10891 , w8891 );
nor ( w10893 , w9012 , w9113 );
not ( w10894 , w10893 );
and ( w10895 , w10894 , w8891 );
and ( w10896 , w10892 , w10895 );
and ( w10897 , w10896 , w8891 );
nor ( w10898 , w10897 , w9027 );
not ( w10899 , w10885 );
and ( w10900 , w10899 , w10898 );
and ( w10901 , w10900 , w9013 );
not ( w10902 , w10901 );
and ( w10903 , w10902 , w9724 );
nor ( w10904 , w10903 , w9249 );
not ( w10905 , w9027 );
and ( w10906 , w10904 , w10905 );
not ( w10907 , w10906 );
and ( w10908 , w10907 , w9122 );
and ( w10909 , w10908 , w8891 );
and ( w10910 , w10909 , w8879 );
and ( w10911 , w10910 , w8891 );
and ( w10912 , w10911 , w11029 );
not ( w10913 , w10912 );
and ( w10914 , w10913 , w8922 );
not ( w10915 , w10914 );
and ( w10916 , w10915 , w9133 );
nor ( w10917 , w10916 , w10871 );
not ( w10918 , w10917 );
and ( w10919 , w10918 , w8891 );
and ( w10920 , w10919 , w10139 );
not ( w10921 , w10920 );
and ( w10922 , w10921 , w8922 );
and ( w10923 , w10922 , w10898 );
not ( w10924 , w9060 );
and ( w10925 , w10924 , w8922 );
nor ( w10926 , w10925 , w10778 );
and ( w10927 , w10926 , w8891 );
nor ( w10928 , w10927 , w8936 );
not ( w10929 , w10928 );
and ( w10930 , w10929 , w8891 );
not ( w10931 , w10930 );
and ( w10932 , w10931 , w8865 );
and ( w10933 , w10987 , w8865 );
and ( w10934 , w10933 , w9069 );
and ( w10935 , w10932 , w10934 );
and ( w10936 , w10935 , w9069 );
not ( w10937 , w10936 );
and ( w10938 , w10937 , w8891 );
nor ( w10939 , w10938 , w8988 );
not ( w10940 , w10939 );
and ( w10941 , w10940 , w8879 );
and ( w10942 , w10941 , w8891 );
nor ( w10943 , w10942 , w8994 );
not ( w10944 , w10943 );
and ( w10945 , w10944 , w8891 );
nor ( w10946 , w10945 , w9012 );
not ( w10947 , w10946 );
and ( w10948 , w10947 , w8891 );
not ( w10949 , w8906 );
and ( w10950 , w10948 , w10949 );
and ( w10951 , w10950 , w8890 );
nor ( w10952 , w10951 , w8909 );
not ( w10953 , w10952 );
and ( w10954 , w10953 , w8891 );
not ( w10955 , w8913 );
and ( w10956 , w10954 , w10955 );
and ( w10957 , w10956 , w8891 );
and ( w10958 , w10957 , w8879 );
and ( w10959 , w10958 , w8891 );
and ( w10960 , w10959 , w11029 );
and ( w10961 , w10960 , w8891 );
and ( w10962 , w10961 , w11078 );
and ( w10963 , w10962 , w9133 );
nor ( w10964 , w10963 , w10871 );
not ( w10965 , w10964 );
and ( w10966 , w10965 , w8891 );
and ( w10967 , w10966 , w10139 );
nor ( w10968 , w8898 , w10967 );
not ( w10969 , w8957 );
and ( w10970 , w10969 , w8977 );
not ( w10971 , w10970 );
and ( w10972 , w10971 , w8865 );
and ( w10973 , w10972 , w10934 );
and ( w10974 , w10973 , w9069 );
and ( w10975 , w10974 , w10301 );
not ( w10976 , w10975 );
and ( w10977 , w10976 , w8891 );
not ( w10978 , w8997 );
and ( w10979 , w10977 , w10978 );
nor ( w10980 , w10979 , w9012 );
not ( w10981 , w10980 );
and ( w10982 , w10981 , w8985 );
and ( w10983 , w10982 , w8891 );
nor ( w10984 , w10983 , w10349 );
nor ( w10985 , w10968 , w10984 );
and ( w10986 , w10985 , w8891 );
not ( w10987 , w9198 );
and ( w10988 , w10987 , w10778 );
not ( w10989 , w10988 );
and ( w10990 , w10989 , w8891 );
not ( w10991 , w10990 );
and ( w10992 , w10991 , w8865 );
and ( w10993 , w10992 , w8933 );
not ( w10994 , w8936 );
and ( w10995 , w10993 , w10994 );
not ( w10996 , w10995 );
and ( w10997 , w10996 , w8879 );
and ( w10998 , w10997 , w8891 );
not ( w10999 , w8989 );
and ( w11000 , w10998 , w10999 );
nor ( w11001 , w11000 , w8994 );
nor ( w11002 , w11001 , w8997 );
nor ( w11003 , w11002 , w8988 );
not ( w11004 , w9012 );
and ( w11005 , w11003 , w11004 );
not ( w11006 , w11005 );
and ( w11007 , w11006 , w8891 );
and ( w11008 , w11007 , w8879 );
and ( w11009 , w11008 , w9113 );
and ( w11010 , w10986 , w11009 );
and ( w11011 , w11010 , w8891 );
and ( w11012 , w11011 , w9113 );
and ( w11013 , w11012 , w8891 );
and ( w11014 , w11013 , w11078 );
and ( w11015 , w11014 , w9133 );
nor ( w11016 , w11015 , w10871 );
not ( w11017 , w11016 );
and ( w11018 , w11017 , w8891 );
and ( w11019 , w11018 , w10139 );
not ( w11020 , w11019 );
and ( w11021 , w10923 , w11020 );
not ( w11022 , w9249 );
and ( w11023 , w11021 , w11022 );
not ( w11024 , w11023 );
and ( w11025 , w11024 , w9122 );
and ( w11026 , w11025 , w8891 );
and ( w11027 , w11026 , w8879 );
and ( w11028 , w11027 , w8891 );
not ( w11029 , w9458 );
and ( w11030 , w11028 , w11029 );
not ( w11031 , w11030 );
and ( w11032 , w11031 , w8922 );
not ( w11033 , w11032 );
and ( w11034 , w11033 , w9133 );
nor ( w11035 , w11034 , w10871 );
not ( w11036 , w11035 );
and ( w11037 , w11036 , w8891 );
and ( w11038 , w11037 , w10139 );
not ( w11039 , w9035 );
and ( w11040 , w11039 , w11038 );
nor ( w11041 , w11040 , w9027 );
not ( w11042 , w11041 );
and ( w11043 , w11042 , w9122 );
not ( w11044 , w11043 );
and ( w11045 , w11044 , w8922 );
not ( w11046 , w10871 );
and ( w11047 , w11045 , w11046 );
not ( w11048 , w9029 );
and ( w11049 , w11048 , w11047 );
and ( w11050 , w11049 , w8922 );
nor ( w11051 , w11050 , w9132 );
and ( w11052 , w11051 , w9133 );
nor ( w11053 , w11052 , w10871 );
not ( w11054 , w11053 );
and ( w11055 , w11054 , w8891 );
and ( w11056 , w11055 , w10139 );
nor ( w11057 , w8924 , w11056 );
not ( w11058 , w11057 );
and ( w11059 , w11058 , w8891 );
and ( w11060 , w11059 , w11078 );
and ( w11061 , w11060 , w9133 );
nor ( w11062 , w11061 , w10871 );
not ( w11063 , w8899 );
and ( w11064 , w11063 , w11062 );
and ( w11065 , w11064 , w9241 );
not ( w11066 , w11065 );
and ( w11067 , w11066 , w8891 );
nor ( w11068 , w11067 , w9249 );
not ( w11069 , w11068 );
and ( w11070 , w11069 , w8891 );
and ( w11071 , w11070 , w8879 );
not ( w11072 , w11071 );
and ( w11073 , w11072 , w9458 );
nor ( w11074 , w11073 , w8923 );
nor ( w11075 , w11074 , w11056 );
not ( w11076 , w11075 );
and ( w11077 , w11076 , w8891 );
not ( w11078 , w9132 );
and ( w11079 , w11077 , w11078 );
and ( w11080 , w11079 , w9133 );
nor ( w11081 , w11080 , w10871 );
and ( t_2 , w8865 , w11081 );
not ( w11082 , w5 );
and ( w11083 , w11082 , g5 );
nor ( w11084 , w11083 , g7 );
and ( w11085 , w3 , g7 );
nor ( w11086 , w11084 , w11085 );
and ( w11087 , w2551 , w11092 );
nor ( w11088 , w11087 , w4179 );
and ( w11089 , w11088 , w12612 );
nor ( w11090 , w11087 , g7 );
nor ( w11091 , w11085 , w11090 );
not ( w11092 , g5 );
and ( w11093 , w11091 , w11092 );
nor ( w11094 , w4 , w11093 );
nor ( w11095 , w11089 , w11094 );
not ( w11096 , w11087 );
and ( w11097 , w11096 , g5 );
not ( w11098 , w11097 );
and ( w11099 , w11098 , g5 );
nor ( w11100 , w11095 , w11099 );
and ( w11101 , w11100 , w12612 );
not ( w11102 , w11086 );
and ( w11103 , w11102 , w11101 );
and ( w11104 , w11103 , w12612 );
and ( w11105 , w13367 , w310 );
and ( w11106 , w3452 , w13536 );
nor ( w11107 , w11085 , w219 );
and ( w11108 , w11107 , w11245 );
and ( w11109 , w11106 , w11108 );
nor ( w11110 , w3456 , w11109 );
nor ( w11111 , w11110 , w11099 );
and ( w11112 , w11111 , w11108 );
not ( w11113 , w11112 );
and ( w11114 , g31 , w11113 );
and ( w11115 , w11105 , w11114 );
and ( w11116 , g8 , w13590 );
and ( w11117 , w11116 , w13536 );
and ( w11118 , w11117 , w12612 );
nor ( w11119 , g9 , w11118 );
and ( w11120 , w12195 , w41 );
nor ( w11121 , w11120 , w48 );
and ( w11122 , w56 , w13536 );
and ( w11123 , w11122 , w12612 );
and ( w11124 , w56 , w11335 );
nor ( w11125 , w11124 , w11099 );
and ( w11126 , w11125 , w12612 );
and ( w11127 , w11126 , w13536 );
and ( w11128 , w11127 , w12612 );
and ( w11129 , w11128 , w13536 );
and ( w11130 , w11129 , w12612 );
nor ( w11131 , w7476 , w274 );
not ( w11132 , w428 );
and ( w11133 , w11131 , w11132 );
nor ( w11134 , w11133 , w272 );
nor ( w11135 , w11134 , w31 );
nor ( w11136 , w11135 , w35 );
nor ( w11137 , w11136 , w37 );
not ( w11138 , w11137 );
and ( w11139 , w11130 , w11138 );
not ( w11140 , w39 );
and ( w11141 , w11139 , w11140 );
and ( w11142 , w11141 , w12117 );
and ( w11143 , w146 , w12950 );
and ( w11144 , w11142 , w12119 );
nor ( w11145 , w11144 , w43 );
and ( w11146 , w11145 , w12142 );
nor ( w11147 , w11146 , w18 );
and ( w11148 , w11094 , w13536 );
and ( w11149 , w11148 , w12612 );
nor ( w11150 , w11147 , w11149 );
nor ( w11151 , w41 , w11099 );
and ( w11152 , w11151 , w12612 );
not ( w11153 , w11150 );
and ( w11154 , w11153 , w11152 );
nor ( w11155 , w105 , w11099 );
and ( w11156 , w11155 , w12612 );
and ( w11157 , w11154 , w11156 );
nor ( w11158 , w11157 , w11094 );
nor ( w11159 , w11158 , w11099 );
nor ( w11160 , w11085 , w11104 );
nor ( w11161 , w11160 , w53 );
nor ( w11162 , w11159 , w11161 );
and ( w11163 , w18 , g12 );
and ( w11164 , w18 , g13 );
nor ( w11165 , w11163 , w11164 );
not ( w11166 , w105 );
and ( w11167 , w11165 , w11166 );
nor ( w11168 , w18 , w105 );
nor ( w11169 , w11167 , w11168 );
and ( w11170 , w11169 , w12057 );
and ( w11171 , w11170 , w12037 );
and ( w11172 , w11171 , w11112 );
nor ( w11173 , w485 , w11099 );
and ( w11174 , w11173 , w11108 );
and ( w11175 , w11172 , w11174 );
and ( w11176 , w377 , w11175 );
nor ( w11177 , w11176 , w11149 );
and ( w11178 , w11177 , w12950 );
nor ( w11179 , w11178 , w11099 );
and ( w11180 , w11179 , w12612 );
nor ( w11181 , w11094 , w11175 );
and ( w11182 , w11169 , w12720 );
and ( w11183 , w11182 , w12057 );
and ( w11184 , w11183 , w11174 );
nor ( w11185 , w1934 , w1853 );
nor ( w11186 , g39 , g13 );
nor ( w11187 , w11185 , w11186 );
nor ( w11188 , w11187 , w11108 );
nor ( w11189 , w11188 , w11099 );
and ( w11190 , w11189 , w13331 );
and ( w11191 , w11190 , g47 );
and ( w11192 , w11191 , w13257 );
and ( w11193 , g48 , g31 );
and ( w11194 , w11192 , w13042 );
and ( w11195 , w11187 , w11094 );
and ( w11196 , w11194 , w11195 );
nor ( w11197 , g36 , g11 );
not ( w11198 , w11197 );
and ( w11199 , w11198 , w11094 );
and ( w11200 , w11196 , w11199 );
nor ( w11201 , w11200 , w11108 );
nor ( w11202 , w11201 , w11099 );
and ( w11203 , w11170 , g32 );
and ( w11204 , w11203 , w11174 );
and ( w11205 , w11204 , w11112 );
nor ( w11206 , w11094 , w11205 );
not ( w11207 , w11206 );
and ( w11208 , w11202 , w11207 );
and ( w11209 , w11208 , g33 );
not ( w11210 , w11185 );
and ( w11211 , w11210 , w11195 );
and ( w11212 , w11211 , w13042 );
and ( w11213 , w11212 , w13257 );
and ( w11214 , w11213 , w11199 );
and ( w11215 , w11214 , w11094 );
and ( w11216 , w11215 , w13331 );
not ( w11217 , g47 );
and ( w11218 , w11216 , w11217 );
not ( w11219 , w11167 );
and ( w11220 , w11219 , w11174 );
and ( w11221 , w11220 , w11112 );
and ( w11222 , w11221 , w11525 );
and ( w11223 , w11222 , w13536 );
and ( w11224 , w11223 , w11108 );
and ( w11225 , w11224 , w12057 );
not ( w11226 , g32 );
and ( w11227 , w11225 , w11226 );
nor ( w11228 , w11218 , w11227 );
nor ( w11229 , w11228 , g33 );
nor ( w11230 , w11209 , w11229 );
not ( w11231 , w11184 );
and ( w11232 , w11231 , w11230 );
nor ( w11233 , w11232 , g29 );
nor ( w11234 , w11094 , w11233 );
and ( w11235 , w11181 , w11234 );
nor ( w11236 , w11235 , g29 );
and ( w11237 , w53 , w11654 );
nor ( w11238 , w11237 , w11099 );
nor ( w11239 , w312 , g30 );
and ( w11240 , w11239 , w13206 );
and ( w11241 , w255 , w11240 );
and ( w11242 , w11240 , g28 );
and ( w11243 , w11242 , g29 );
nor ( w11244 , w11241 , w11243 );
not ( w11245 , w4179 );
and ( w11246 , w3 , w11245 );
and ( w11247 , w11246 , g5 );
nor ( w11248 , w11247 , w11085 );
not ( w11249 , w11248 );
and ( w11250 , w11249 , w11108 );
nor ( w11251 , w11094 , w11250 );
not ( w11252 , w11085 );
and ( w11253 , w11251 , w11252 );
not ( w11254 , w11253 );
and ( w11255 , w11254 , w11108 );
not ( w11256 , w11255 );
and ( w11257 , w11244 , w11256 );
and ( w11258 , w11525 , w11108 );
not ( w11259 , w11257 );
and ( w11260 , w11259 , w11258 );
not ( w11261 , g10 );
and ( w11262 , w11260 , w11261 );
and ( w11263 , w11262 , w11108 );
and ( w11264 , w11263 , w13477 );
nor ( w11265 , w11094 , w11264 );
not ( w11266 , w11265 );
and ( w11267 , w11238 , w11266 );
nor ( w11268 , w11236 , w11267 );
not ( w11269 , w11180 );
and ( w11270 , w11269 , w11268 );
and ( w11271 , w11270 , w11585 );
nor ( w11272 , w11271 , w11099 );
and ( w11273 , w11272 , w12612 );
and ( w11274 , w11162 , w12930 );
nor ( w11275 , w11274 , w53 );
not ( w11276 , w11275 );
and ( w11277 , w11121 , w11276 );
and ( w11278 , w255 , w12612 );
nor ( w11279 , w5 , g7 );
nor ( w11280 , w11279 , w222 );
and ( w11281 , w11280 , w13536 );
and ( w11282 , w11281 , w11094 );
and ( w11283 , w13536 , w11255 );
and ( w11284 , w11283 , w11108 );
nor ( w11285 , w11282 , w11284 );
not ( w11286 , w11278 );
and ( w11287 , w11286 , w11285 );
nor ( w11288 , w19 , w11287 );
nor ( w11289 , w11149 , w11094 );
nor ( w11290 , w11289 , w11099 );
and ( w11291 , w11290 , w12612 );
nor ( w11292 , w11149 , w11291 );
and ( w11293 , w11292 , w12950 );
nor ( w11294 , w11293 , w11099 );
and ( w11295 , w11294 , w12612 );
not ( w11296 , w11295 );
and ( w11297 , w11292 , w11296 );
and ( w11298 , w11297 , w12950 );
nor ( w11299 , w11298 , w11099 );
and ( w11300 , w11299 , w12612 );
and ( w11301 , w11292 , w11671 );
and ( w11302 , w11301 , w12725 );
and ( w11303 , w11302 , w12950 );
nor ( w11304 , w11303 , w11099 );
and ( w11305 , w11304 , w12612 );
nor ( w11306 , w11305 , w11149 );
and ( w11307 , w11306 , w12950 );
nor ( w11308 , w11307 , w11099 );
and ( w11309 , w11308 , w12612 );
nor ( w11310 , w11149 , w11309 );
and ( w11311 , g10 , w12720 );
and ( w11312 , w11311 , g11 );
and ( w11313 , w11312 , w11533 );
and ( w11314 , w11313 , w11797 );
and ( w11315 , w12720 , g10 );
and ( w11316 , w11315 , g11 );
and ( w11317 , w11316 , w11533 );
and ( w11318 , w11317 , w11797 );
and ( w11319 , w11318 , w11156 );
not ( w11320 , w11319 );
and ( w11321 , w11320 , w11268 );
and ( w11322 , w11321 , w12950 );
nor ( w11323 , w11322 , w11099 );
and ( w11324 , w11323 , w12612 );
nor ( w11325 , w11314 , w11324 );
nor ( w11326 , w20 , w11119 );
and ( w11327 , w21 , w13536 );
and ( w11328 , w11327 , w12612 );
nor ( w11329 , w428 , w11099 );
and ( w11330 , w11329 , w12612 );
and ( w11331 , w11328 , w11330 );
and ( w11332 , w272 , w13536 );
and ( w11333 , w11332 , w12612 );
nor ( w11334 , w11331 , w11333 );
not ( w11335 , w11123 );
and ( w11336 , w11334 , w11335 );
nor ( w11337 , w31 , w11099 );
and ( w11338 , w11337 , w12612 );
not ( w11339 , w11336 );
and ( w11340 , w11339 , w11338 );
nor ( w11341 , w274 , w11099 );
and ( w11342 , w11341 , w12612 );
and ( w11343 , w11340 , w11342 );
and ( w11344 , w35 , w13536 );
and ( w11345 , w11344 , w12612 );
nor ( w11346 , w11343 , w11345 );
not ( w11347 , w33 );
and ( w11348 , w11347 , w11346 );
nor ( w11349 , w37 , w11099 );
and ( w11350 , w11349 , w12612 );
not ( w11351 , w11348 );
and ( w11352 , w11351 , w11350 );
and ( w11353 , w11352 , w13536 );
and ( w11354 , w11353 , w12612 );
and ( w11355 , w39 , w13536 );
and ( w11356 , w11355 , w12612 );
nor ( w11357 , w11354 , w11356 );
not ( w11358 , w11357 );
and ( w11359 , w11358 , w11152 );
and ( w11360 , w45 , w13536 );
and ( w11361 , w11360 , w12612 );
nor ( w11362 , w11359 , w11361 );
and ( w11363 , w11326 , w11515 );
and ( w11364 , w11363 , w12720 );
nor ( w11365 , w43 , w11099 );
and ( w11366 , w11365 , w12612 );
and ( w11367 , w11364 , w11366 );
nor ( w11368 , w11367 , w11149 );
not ( w11369 , w11368 );
and ( w11370 , w11369 , w377 );
nor ( w11371 , w11370 , w11149 );
and ( w11372 , w11306 , w11268 );
and ( w11373 , w11372 , w12725 );
nor ( w11374 , w11373 , w11099 );
and ( w11375 , w11374 , w12612 );
nor ( w11376 , w11375 , w11305 );
and ( w11377 , w11376 , w12725 );
and ( w11378 , w11377 , w11268 );
and ( w11379 , w11378 , w12725 );
and ( w11380 , w11379 , w12950 );
nor ( w11381 , w11380 , w11099 );
and ( w11382 , w11381 , w12612 );
nor ( w11383 , w11382 , w11305 );
and ( w11384 , w11383 , w12725 );
and ( w11385 , w11384 , w11268 );
and ( w11386 , w11385 , w12950 );
nor ( w11387 , w11386 , w11099 );
and ( w11388 , w11387 , w12612 );
not ( w11389 , w11388 );
and ( w11390 , w11306 , w11389 );
and ( w11391 , w11390 , w12725 );
and ( w11392 , w12725 , w11268 );
and ( w11393 , w11392 , w12950 );
nor ( w11394 , w11393 , w11099 );
and ( w11395 , w11394 , w12612 );
not ( w11396 , w11395 );
and ( w11397 , w11391 , w11396 );
and ( w11398 , w11397 , w11268 );
and ( w11399 , w11398 , w12950 );
nor ( w11400 , w11399 , w11099 );
nor ( w11401 , w11400 , w11149 );
nor ( w11402 , w11401 , w53 );
and ( w11403 , w11371 , w11420 );
not ( w11404 , w11403 );
and ( w11405 , w11404 , w11156 );
not ( w11406 , w11405 );
and ( w11407 , w11406 , w11268 );
and ( w11408 , w11407 , w12950 );
nor ( w11409 , w11408 , w11099 );
nor ( w11410 , w11409 , w11149 );
and ( w11411 , w11173 , w12612 );
not ( w11412 , w11410 );
and ( w11413 , w11412 , w11411 );
and ( w11414 , w11413 , w12612 );
not ( w11415 , w11414 );
and ( w11416 , w11325 , w11415 );
not ( w11417 , w11416 );
and ( w11418 , w11417 , w377 );
nor ( w11419 , w11418 , w11149 );
not ( w11420 , w11402 );
and ( w11421 , w11419 , w11420 );
not ( w11422 , w11421 );
and ( w11423 , w11422 , w11156 );
not ( w11424 , w11423 );
and ( w11425 , w11424 , w11268 );
and ( w11426 , w11425 , w12950 );
nor ( w11427 , w11426 , w11099 );
and ( w11428 , w11427 , w12612 );
not ( w11429 , w11428 );
and ( w11430 , w11310 , w11429 );
and ( w11431 , w11430 , w11268 );
and ( w11432 , w11431 , w12950 );
nor ( w11433 , w11432 , w11099 );
and ( w11434 , w11433 , w12612 );
nor ( w11435 , w11149 , w11434 );
and ( w11436 , w11326 , w377 );
nor ( w11437 , w11436 , w11149 );
nor ( w11438 , w11437 , w11362 );
and ( w11439 , w11438 , w11366 );
nor ( w11440 , w11439 , w11149 );
not ( w11441 , w11440 );
and ( w11442 , w11441 , w11156 );
nor ( w11443 , w11442 , w11094 );
nor ( w11444 , w11443 , w11099 );
nor ( w11445 , w11444 , w11149 );
not ( w11446 , w11445 );
and ( w11447 , w11446 , w11411 );
and ( w11448 , w11447 , w12612 );
nor ( w11449 , w11448 , w11309 );
nor ( w11450 , w377 , w11149 );
not ( w11451 , w11450 );
and ( w11452 , w11451 , g10 );
and ( w11453 , w11452 , g11 );
and ( w11454 , w11453 , w11533 );
and ( w11455 , w11454 , w11797 );
nor ( w11456 , w11455 , w11094 );
nor ( w11457 , w11456 , w11099 );
and ( w11458 , w11457 , w12612 );
not ( w11459 , w11458 );
and ( w11460 , w11449 , w11459 );
not ( w11461 , w11460 );
and ( w11462 , w11461 , w11156 );
nor ( w11463 , w11462 , w11180 );
nor ( w11464 , w11463 , w11114 );
nor ( w11465 , w11464 , w11434 );
and ( w11466 , w11465 , w12950 );
nor ( w11467 , w11466 , w11099 );
nor ( w11468 , w11467 , w11149 );
and ( w11469 , w11292 , w11671 );
and ( w11470 , w11469 , w11114 );
nor ( w11471 , w11114 , g28 );
and ( w11472 , w11471 , w13333 );
and ( w11473 , w11472 , w12037 );
and ( w11474 , w11473 , w11174 );
nor ( w11475 , w11474 , w11236 );
and ( w11476 , w11475 , w11585 );
and ( w11477 , w11476 , g8 );
and ( w11478 , w11477 , g9 );
and ( w11479 , w11478 , w12950 );
nor ( w11480 , w11168 , w11479 );
and ( w11481 , w11480 , g8 );
and ( w11482 , w11481 , g9 );
nor ( w11483 , w11482 , w11094 );
nor ( w11484 , w11483 , w11099 );
and ( w11485 , w11484 , w12612 );
not ( w11486 , w11485 );
and ( w11487 , w11470 , w11486 );
not ( w11488 , w11487 );
and ( w11489 , w11488 , g13 );
nor ( w11490 , w11489 , g12 );
and ( w11491 , w11490 , w12725 );
and ( w11492 , w11301 , w11114 );
nor ( w11493 , w11492 , w11119 );
and ( w11494 , w11493 , w11515 );
nor ( w11495 , w11494 , w11149 );
not ( w11496 , w11495 );
and ( w11497 , w11496 , w11366 );
nor ( w11498 , w11497 , w11485 );
and ( w11499 , w11498 , w12725 );
not ( w11500 , w11499 );
and ( w11501 , w11500 , w377 );
and ( w11502 , w11501 , w11411 );
not ( w11503 , w11502 );
and ( w11504 , w11503 , g12 );
not ( w11505 , w11504 );
and ( w11506 , w11505 , w11156 );
nor ( w11507 , w11506 , w11094 );
nor ( w11508 , w11507 , w11099 );
and ( w11509 , w11508 , w12612 );
not ( w11510 , w11491 );
and ( w11511 , w11510 , w11509 );
not ( w11512 , w11511 );
and ( w11513 , w11512 , w11268 );
and ( w11514 , w11513 , w11114 );
not ( w11515 , w11362 );
and ( w11516 , w11515 , w11366 );
nor ( w11517 , w11516 , w11485 );
nor ( w11518 , w11517 , w11119 );
and ( w11519 , w11518 , g13 );
nor ( w11520 , w11519 , g12 );
not ( w11521 , w11520 );
and ( w11522 , w11521 , w11411 );
and ( w11523 , w11522 , w11509 );
and ( w11524 , w11523 , w11156 );
not ( w11525 , w11168 );
and ( w11526 , w11174 , w11525 );
nor ( w11527 , w11526 , w11267 );
not ( w11528 , w11527 );
and ( w11529 , w11528 , w105 );
nor ( w11530 , w11529 , w11094 );
not ( w11531 , w11524 );
and ( w11532 , w11531 , w11530 );
not ( w11533 , g12 );
and ( w11534 , w11114 , w11533 );
and ( w11535 , w11534 , w11797 );
and ( w11536 , w11797 , w11509 );
not ( w11537 , w11535 );
and ( w11538 , w11537 , w11536 );
and ( w11539 , w11538 , w11509 );
not ( w11540 , w11539 );
and ( w11541 , w11540 , w11268 );
and ( w11542 , w11541 , w11114 );
nor ( w11543 , w19 , g12 );
and ( w11544 , w11543 , w11797 );
not ( w11545 , w11544 );
and ( w11546 , w11545 , w11536 );
and ( w11547 , w11546 , w11509 );
and ( w11548 , w11547 , w11156 );
and ( w11549 , w11548 , w377 );
and ( w11550 , w11549 , w13536 );
and ( w11551 , w11550 , w12612 );
and ( w11552 , w11551 , w11536 );
not ( w11553 , w11552 );
and ( w11554 , w11553 , w11530 );
not ( w11555 , w11554 );
and ( w11556 , w11555 , w377 );
nor ( w11557 , w11556 , w11094 );
nor ( w11558 , w11557 , w11099 );
and ( w11559 , w11558 , w12612 );
not ( w11560 , w11542 );
and ( w11561 , w11560 , w11559 );
nor ( w11562 , w11561 , w11094 );
nor ( w11563 , w11562 , w11099 );
and ( w11564 , w11563 , w12612 );
and ( w11565 , w11532 , w11574 );
not ( w11566 , w11565 );
and ( w11567 , w11566 , w377 );
nor ( w11568 , w11567 , w11094 );
nor ( w11569 , w11568 , w11099 );
and ( w11570 , w11569 , w12612 );
not ( w11571 , w11514 );
and ( w11572 , w11571 , w11570 );
nor ( w11573 , w11572 , w11149 );
not ( w11574 , w11564 );
and ( w11575 , w11573 , w11574 );
and ( w11576 , w11575 , w12950 );
nor ( w11577 , w11576 , w11099 );
and ( w11578 , w11577 , w12612 );
nor ( w11579 , w11149 , w11578 );
and ( w11580 , w11579 , w12950 );
nor ( w11581 , w11580 , w11099 );
and ( w11582 , w11581 , w12612 );
and ( w11583 , w11306 , w11595 );
and ( w11584 , w11450 , w11268 );
not ( w11585 , w11267 );
and ( w11586 , w11584 , w11585 );
nor ( w11587 , w11586 , w11530 );
and ( w11588 , w11587 , w13536 );
and ( w11589 , w11588 , w12612 );
not ( w11590 , w11589 );
and ( w11591 , w11583 , w11590 );
nor ( w11592 , w11591 , w11114 );
nor ( w11593 , w11388 , w11305 );
and ( w11594 , w11593 , w12725 );
not ( w11595 , w11582 );
and ( w11596 , w11594 , w11595 );
and ( w11597 , w11596 , w11268 );
and ( w11598 , w11597 , w12725 );
and ( w11599 , w11598 , w11605 );
and ( w11600 , w11599 , w12950 );
nor ( w11601 , w11600 , w11099 );
and ( w11602 , w11601 , w12612 );
nor ( w11603 , w11592 , w11602 );
and ( w11604 , w11603 , w12725 );
not ( w11605 , w11578 );
and ( w11606 , w11604 , w11605 );
and ( w11607 , w11606 , w12950 );
nor ( w11608 , w11607 , w11099 );
and ( w11609 , w11608 , w12612 );
not ( w11610 , w11609 );
and ( w11611 , w11468 , w11610 );
nor ( w11612 , w11611 , w53 );
and ( w11613 , w11435 , w11818 );
and ( w11614 , w11619 , w11613 );
and ( w11615 , w11614 , w11818 );
nor ( w11616 , w11615 , w53 );
not ( w11617 , w11616 );
and ( w11618 , w11617 , w11285 );
not ( w11619 , w11288 );
and ( w11620 , w11619 , w11618 );
and ( w11621 , w11620 , w11818 );
and ( w11622 , w11621 , w12950 );
nor ( w11623 , w11622 , w11099 );
and ( w11624 , w11623 , w12612 );
not ( w11625 , w11624 );
and ( w11626 , w11625 , w11285 );
and ( w11627 , w11277 , w11626 );
not ( w11628 , w11627 );
and ( w11629 , w11628 , w11174 );
and ( w11630 , w12725 , w11285 );
not ( w11631 , w11629 );
and ( w11632 , w11631 , w11630 );
not ( w11633 , w11632 );
and ( w11634 , w11633 , w11156 );
and ( w11635 , w19 , w12612 );
not ( w11636 , w11635 );
and ( w11637 , w11636 , w11285 );
not ( w11638 , w11637 );
and ( w11639 , w11634 , w11638 );
nor ( w11640 , w11639 , w11094 );
nor ( w11641 , w11161 , w11273 );
and ( w11642 , w11641 , w12950 );
nor ( w11643 , w11642 , w11099 );
and ( w11644 , w11643 , w12612 );
nor ( w11645 , w11644 , w11161 );
and ( w11646 , w11645 , w12725 );
and ( w11647 , w11646 , w11829 );
and ( w11648 , w11647 , w12947 );
and ( w11649 , w11648 , w12930 );
and ( w11650 , w11649 , w12950 );
nor ( w11651 , w11650 , w11099 );
and ( w11652 , w11651 , w12612 );
and ( w11653 , g47 , g33 );
not ( w11654 , w11108 );
and ( w11655 , w11653 , w11654 );
nor ( w11656 , w11655 , w11099 );
and ( w11657 , w13042 , w11656 );
nor ( w11658 , w11230 , g29 );
nor ( w11659 , w11657 , w11658 );
nor ( w11660 , w11659 , g45 );
and ( w11661 , w11660 , w13257 );
and ( w11662 , w11661 , w11195 );
and ( w11663 , w11662 , w11199 );
nor ( w11664 , w11663 , w11108 );
not ( w11665 , w11664 );
and ( w11666 , w11665 , w11189 );
and ( w11667 , w11666 , w13536 );
and ( w11668 , w11667 , w11236 );
and ( w11669 , w11668 , w13333 );
nor ( w11670 , w11669 , w11267 );
not ( w11671 , w11300 );
and ( w11672 , w11671 , w11670 );
and ( w11673 , w11672 , w12725 );
and ( w11674 , w11673 , w12947 );
and ( w11675 , w11674 , w12725 );
and ( w11676 , w11675 , w11829 );
and ( w11677 , w11676 , w12947 );
and ( w11678 , w11677 , w12930 );
and ( w11679 , w11674 , w11678 );
and ( w11680 , w11679 , w12725 );
and ( w11681 , w11680 , w11829 );
and ( w11682 , w11681 , w12947 );
and ( w11683 , w11682 , w12930 );
nor ( w11684 , w11161 , w11149 );
and ( w11685 , w11684 , w12950 );
nor ( w11686 , w11685 , w11099 );
nor ( w11687 , w11686 , w11644 );
and ( w11688 , w11687 , w12947 );
and ( w11689 , w11688 , w12930 );
nor ( w11690 , w11689 , w53 );
nor ( w11691 , w11690 , w11161 );
and ( w11692 , w11691 , w12725 );
and ( w11693 , w11692 , w12950 );
nor ( w11694 , w11693 , w11099 );
nor ( w11695 , w11694 , w11644 );
and ( w11696 , w11695 , w12947 );
and ( w11697 , w11696 , w12930 );
nor ( w11698 , w11697 , w53 );
and ( w11699 , w11683 , w11883 );
and ( w11700 , w11699 , w11678 );
and ( w11701 , w11700 , w12725 );
nor ( w11702 , w11149 , w11652 );
and ( w11703 , g36 , g11 );
and ( w11704 , w11703 , w11795 );
and ( w11705 , w11704 , w11797 );
nor ( w11706 , g42 , g21 );
nor ( w11707 , g40 , g17 );
not ( w11708 , w11707 );
and ( w11709 , w11708 , g41 );
and ( w11710 , w11709 , g15 );
and ( w11711 , g37 , g19 );
and ( w11712 , w11711 , w11094 );
nor ( w11713 , w11712 , w11284 );
not ( w11714 , w11710 );
and ( w11715 , w11714 , w11713 );
and ( w11716 , g40 , g17 );
and ( w11717 , w11716 , w11094 );
nor ( w11718 , w11717 , w11284 );
and ( w11719 , w11715 , w11718 );
nor ( w11720 , g37 , g19 );
and ( w11721 , w13013 , w11094 );
nor ( w11722 , w11721 , w11284 );
nor ( w11723 , w11719 , w11722 );
and ( w11724 , w11723 , w11094 );
nor ( w11725 , w11724 , w11284 );
nor ( w11726 , w11706 , w11725 );
nor ( w11727 , w11726 , w11284 );
and ( w11728 , g42 , g21 );
and ( w11729 , w11728 , w11094 );
not ( w11730 , w11729 );
and ( w11731 , w11727 , w11730 );
not ( w11732 , w9084 );
and ( w11733 , w11732 , w11094 );
nor ( w11734 , w11733 , w11284 );
nor ( w11735 , w11731 , w11734 );
nor ( w11736 , w11735 , w11284 );
and ( w11737 , w9213 , w11094 );
not ( w11738 , w11737 );
and ( w11739 , w11736 , w11738 );
and ( w11740 , w11741 , g25 );
not ( w11741 , w11739 );
and ( w11742 , w11741 , g38 );
and ( w11743 , w11742 , w11094 );
nor ( w11744 , w11743 , w11284 );
not ( w11745 , w11740 );
and ( w11746 , w11745 , w11744 );
and ( w11747 , w8983 , w11094 );
and ( w11748 , w11746 , w13503 );
not ( w11749 , w11748 );
and ( w11750 , w11749 , w11094 );
nor ( w11751 , w11750 , w11284 );
and ( w11752 , g44 , g27 );
and ( w11753 , w11752 , w11094 );
not ( w11754 , w11753 );
and ( w11755 , w11751 , w11754 );
and ( w11756 , w11755 , w13584 );
and ( w11757 , w13528 , w11094 );
nor ( w11758 , w11757 , w11284 );
nor ( w11759 , w11756 , w11758 );
not ( w11760 , w1878 );
and ( w11761 , w11760 , w11094 );
nor ( w11762 , w11761 , w11284 );
and ( w11763 , w11759 , w11789 );
nor ( w11764 , w11763 , w11284 );
and ( w11765 , w11189 , w11195 );
and ( w11766 , w11765 , w11094 );
not ( w11767 , w11766 );
and ( w11768 , w11764 , w11767 );
nor ( w11769 , w11768 , w11186 );
and ( w11770 , w11769 , w11199 );
nor ( w11771 , w11770 , w11284 );
not ( w11772 , w11771 );
and ( w11773 , w11772 , w11094 );
nor ( w11774 , w11773 , w11284 );
not ( w11775 , w11705 );
and ( w11776 , w11775 , w11774 );
nor ( w11777 , w11776 , g45 );
and ( w11778 , w11777 , w13333 );
nor ( w11779 , w11778 , w11284 );
nor ( w11780 , w11779 , w11193 );
and ( w11781 , w11780 , w11656 );
nor ( w11782 , w11193 , g45 );
and ( w11783 , w11782 , w13333 );
not ( w11784 , w11783 );
and ( w11785 , w11784 , w11670 );
nor ( w11786 , w11785 , w11756 );
not ( w11787 , w11758 );
and ( w11788 , w11786 , w11787 );
not ( w11789 , w11762 );
and ( w11790 , w11788 , w11789 );
nor ( w11791 , w11790 , w11284 );
nor ( w11792 , w11791 , w11186 );
and ( w11793 , w11783 , g36 );
and ( w11794 , w11793 , g11 );
not ( w11795 , g39 );
and ( w11796 , w11794 , w11795 );
not ( w11797 , g13 );
and ( w11798 , w11796 , w11797 );
not ( w11799 , w11798 );
and ( w11800 , w11799 , w11670 );
not ( w11801 , w11800 );
and ( w11802 , w11801 , w11094 );
nor ( w11803 , w11802 , w11284 );
not ( w11804 , w11792 );
and ( w11805 , w11804 , w11803 );
and ( w11806 , w11805 , w11670 );
not ( w11807 , w11806 );
and ( w11808 , w11807 , w11199 );
nor ( w11809 , w11808 , w11284 );
not ( w11810 , w11809 );
and ( w11811 , w11810 , w11094 );
nor ( w11812 , w11811 , w11284 );
not ( w11813 , w11781 );
and ( w11814 , w11813 , w11812 );
not ( w11815 , w11814 );
and ( w11816 , w11815 , w11094 );
nor ( w11817 , w11816 , w11284 );
not ( w11818 , w11612 );
and ( w11819 , w11817 , w11818 );
and ( w11820 , w11702 , w11819 );
and ( w11821 , w11820 , w12950 );
nor ( w11822 , w11821 , w11099 );
nor ( w11823 , w11822 , w11161 );
and ( w11824 , w11823 , w12930 );
nor ( w11825 , w11824 , w53 );
nor ( w11826 , w11825 , w11161 );
and ( w11827 , w11826 , w11915 );
and ( w11828 , w11827 , w11819 );
not ( w11829 , w11644 );
and ( w11830 , w11828 , w11829 );
and ( w11831 , w11830 , w12947 );
and ( w11832 , w11701 , w11831 );
and ( w11833 , w11832 , w12950 );
nor ( w11834 , w11833 , w11099 );
nor ( w11835 , w11834 , w11161 );
and ( w11836 , w11835 , w12930 );
nor ( w11837 , w11836 , w53 );
nor ( w11838 , w11652 , w11837 );
and ( w11839 , w11838 , w11917 );
and ( w11840 , w12947 , w11285 );
and ( w11841 , w11839 , w11840 );
nor ( w11842 , w312 , w11841 );
and ( w11843 , w11630 , w12950 );
nor ( w11844 , w11843 , w11099 );
and ( w11845 , w11844 , w12612 );
not ( w11846 , w11845 );
and ( w11847 , w11846 , w11285 );
not ( w11848 , w11842 );
and ( w11849 , w11848 , w11847 );
nor ( w11850 , w11652 , w11161 );
and ( w11851 , w11850 , w11285 );
not ( w11852 , w384 );
and ( w11853 , w11852 , w11851 );
and ( w11854 , w11853 , w11850 );
nor ( w11855 , w11854 , w11099 );
and ( w11856 , w11855 , w12612 );
not ( w11857 , w11856 );
and ( w11858 , w11857 , w11285 );
and ( w11859 , w11915 , w11858 );
and ( w11860 , w11859 , w12947 );
and ( w11861 , w11860 , w11285 );
and ( w11862 , w11915 , w11840 );
and ( w11863 , w11862 , w11850 );
and ( w11864 , w11863 , w11915 );
and ( w11865 , w11864 , w11883 );
and ( w11866 , w11917 , w11613 );
nor ( w11867 , w11434 , w11094 );
nor ( w11868 , w11867 , w11099 );
and ( w11869 , w11868 , w12612 );
nor ( w11870 , w11434 , w11869 );
and ( w11871 , w11870 , w12950 );
nor ( w11872 , w11871 , w11099 );
and ( w11873 , w11872 , w12612 );
not ( w11874 , w11873 );
and ( w11875 , w11874 , w11285 );
and ( w11876 , w11866 , w11875 );
and ( w11877 , w11876 , w11285 );
and ( w11878 , w11865 , w11877 );
and ( w11879 , w11878 , w310 );
and ( w11880 , w11879 , w11114 );
and ( w11881 , w11858 , w11840 );
and ( w11882 , w11881 , w11915 );
not ( w11883 , w11698 );
and ( w11884 , w11882 , w11883 );
and ( w11885 , w11460 , w11917 );
and ( w11886 , w11885 , w11613 );
and ( w11887 , w11870 , g30 );
nor ( w11888 , w11887 , g31 );
nor ( w11889 , w11888 , w11094 );
nor ( w11890 , w11889 , w11099 );
and ( w11891 , w11890 , w12612 );
not ( w11892 , w11891 );
and ( w11893 , w11892 , w11285 );
and ( w11894 , w11870 , w11893 );
and ( w11895 , w11894 , w12950 );
nor ( w11896 , w11895 , w11099 );
and ( w11897 , w11896 , w12612 );
not ( w11898 , w11897 );
and ( w11899 , w11898 , w11285 );
and ( w11900 , w11886 , w11899 );
and ( w11901 , w310 , w12612 );
not ( w11902 , w11901 );
and ( w11903 , w11902 , w11285 );
and ( w11904 , w11900 , w11903 );
not ( w11905 , w11904 );
and ( w11906 , w11905 , w11156 );
nor ( w11907 , w11906 , w11094 );
nor ( w11908 , w11907 , w11099 );
nor ( w11909 , w11908 , w11273 );
nor ( w11910 , w11909 , w53 );
not ( w11911 , w11910 );
and ( w11912 , w11911 , w11285 );
and ( w11913 , w11884 , w11912 );
and ( w11914 , w11913 , w11903 );
not ( w11915 , w11652 );
and ( w11916 , w11700 , w11915 );
not ( w11917 , w11434 );
and ( w11918 , w11916 , w11917 );
and ( w11919 , w11918 , w12725 );
and ( w11920 , w11918 , w12529 );
nor ( w11921 , w384 , w53 );
not ( w11922 , w11921 );
and ( w11923 , w11922 , w11285 );
and ( w11924 , w11920 , w11923 );
and ( w11925 , w11924 , w12725 );
nor ( w11926 , w11925 , w11287 );
not ( w11927 , w11926 );
and ( w11928 , w11927 , w11831 );
and ( w11929 , w11928 , w12950 );
nor ( w11930 , w11929 , w11099 );
nor ( w11931 , w11930 , w11161 );
and ( w11932 , w11931 , w12930 );
nor ( w11933 , w11932 , w53 );
not ( w11934 , w11933 );
and ( w11935 , w11934 , w11285 );
and ( w11936 , w11919 , w11935 );
and ( w11937 , w11936 , w12529 );
and ( w11938 , w11937 , w12199 );
and ( w11939 , w11938 , w13206 );
and ( w11940 , w11939 , w12725 );
and ( w11941 , w11940 , w11831 );
and ( w11942 , w11941 , w12950 );
nor ( w11943 , w11942 , w11099 );
nor ( w11944 , w11943 , w11161 );
and ( w11945 , w11944 , w12930 );
nor ( w11946 , w11945 , w53 );
not ( w11947 , w11946 );
and ( w11948 , w11947 , w11285 );
nor ( w11949 , w11914 , w11948 );
not ( w11950 , w11949 );
and ( w11951 , w11950 , w11831 );
nor ( w11952 , w11951 , w11099 );
nor ( w11953 , w11952 , w11161 );
nor ( w11954 , w11953 , w53 );
not ( w11955 , w11954 );
and ( w11956 , w11955 , w11285 );
nor ( w11957 , w11880 , w11956 );
not ( w11958 , w11957 );
and ( w11959 , w11958 , w11831 );
and ( w11960 , w11959 , w12950 );
nor ( w11961 , w11960 , w11099 );
nor ( w11962 , w11961 , w11161 );
nor ( w11963 , w11962 , w53 );
not ( w11964 , w11963 );
and ( w11965 , w11964 , w11285 );
and ( w11966 , w11683 , w11965 );
and ( w11967 , w11966 , w11678 );
and ( w11968 , w11877 , w310 );
and ( w11969 , w11968 , w11114 );
nor ( w11970 , w11969 , w11912 );
nor ( w11971 , w11970 , w11094 );
nor ( w11972 , w11971 , w11099 );
and ( w11973 , w11972 , w12612 );
not ( w11974 , w11973 );
and ( w11975 , w11974 , w11285 );
and ( w11976 , w11967 , w11975 );
nor ( w11977 , w11976 , w11948 );
nor ( w11978 , w11977 , w11149 );
and ( w11979 , w11978 , w11831 );
and ( w11980 , w11979 , w12950 );
nor ( w11981 , w11980 , w11099 );
nor ( w11982 , w11981 , w11161 );
and ( w11983 , w11982 , w12930 );
nor ( w11984 , w11983 , w53 );
not ( w11985 , w11984 );
and ( w11986 , w11985 , w11285 );
and ( w11987 , w11861 , w11986 );
and ( w11988 , w11987 , w11840 );
and ( w11989 , w11988 , w11975 );
nor ( w11990 , w11989 , w11948 );
not ( w11991 , w11990 );
and ( w11992 , w11991 , w11831 );
and ( w11993 , w11992 , w12950 );
nor ( w11994 , w11993 , w11099 );
nor ( w11995 , w11994 , w11161 );
nor ( w11996 , w11995 , w53 );
not ( w11997 , w11996 );
and ( w11998 , w11997 , w11285 );
and ( w11999 , w11987 , w11998 );
and ( w12000 , w11999 , w11975 );
nor ( w12001 , w12000 , w11948 );
not ( w12002 , w12001 );
and ( w12003 , w12002 , w11831 );
and ( w12004 , w12003 , w12950 );
nor ( w12005 , w12004 , w11099 );
nor ( w12006 , w12005 , w11161 );
nor ( w12007 , w12006 , w53 );
not ( w12008 , w12007 );
and ( w12009 , w12008 , w11285 );
and ( w12010 , w11849 , w12009 );
and ( w12011 , w12010 , w12725 );
and ( w12012 , w12011 , w11831 );
and ( w12013 , w12012 , w12950 );
nor ( w12014 , w12013 , w11099 );
nor ( w12015 , w12014 , w11161 );
nor ( w12016 , w12015 , w53 );
not ( w12017 , w12016 );
and ( w12018 , w12017 , w11285 );
and ( w12019 , w11640 , w12018 );
nor ( w12020 , w12019 , w11099 );
nor ( w12021 , w12020 , w11104 );
and ( w12022 , w12021 , w12930 );
nor ( w12023 , w12022 , w53 );
not ( w12024 , w11115 );
and ( w12025 , w12024 , w12023 );
and ( w12026 , w12025 , w12562 );
and ( w12027 , w12026 , w377 );
and ( w12028 , w12027 , w12057 );
and ( w12029 , w12028 , w13333 );
nor ( w12030 , w11366 , w43 );
nor ( w12031 , w12030 , w11119 );
nor ( w12032 , w12031 , w48 );
not ( w12033 , w12032 );
and ( w12034 , w12033 , w308 );
and ( w12035 , w12034 , w12717 );
and ( w12036 , w12035 , w308 );
not ( w12037 , w312 );
and ( w12038 , w12037 , w11923 );
not ( w12039 , w12038 );
and ( w12040 , w12039 , g10 );
and ( w12041 , w12040 , g11 );
not ( w12042 , w12041 );
and ( w12043 , w12042 , w11935 );
and ( w12044 , w12043 , w12947 );
nor ( w12045 , w12044 , w53 );
not ( w12046 , w12045 );
and ( w12047 , w12046 , w11285 );
and ( w12048 , w12117 , w41 );
and ( w12049 , w312 , w12612 );
not ( w12050 , w12049 );
and ( w12051 , w12050 , w11285 );
and ( w12052 , w7791 , w12051 );
not ( w12053 , w12052 );
and ( w12054 , w12053 , w11130 );
and ( w12055 , w12054 , w12195 );
and ( w12056 , w12055 , w377 );
not ( w12057 , g28 );
and ( w12058 , w312 , w12057 );
not ( w12059 , w12058 );
and ( w12060 , w12059 , w11923 );
nor ( w12061 , w377 , w53 );
not ( w12062 , w12061 );
and ( w12063 , w12062 , w11285 );
nor ( w12064 , w12060 , w12063 );
and ( w12065 , w12064 , g29 );
nor ( w12066 , w12038 , w12063 );
and ( w12067 , w12066 , g28 );
and ( w12068 , w12067 , w13333 );
and ( w12069 , w12068 , w13536 );
and ( w12070 , w12069 , w12612 );
not ( w12071 , w12070 );
and ( w12072 , w12071 , w11285 );
not ( w12073 , w12065 );
and ( w12074 , w12073 , w12072 );
nor ( w12075 , w12074 , w11099 );
nor ( w12076 , w12075 , w11161 );
nor ( w12077 , w12076 , w53 );
not ( w12078 , w12077 );
and ( w12079 , w12078 , w11285 );
not ( w12080 , w255 );
and ( w12081 , w12080 , w12079 );
and ( w12082 , w12081 , w12072 );
nor ( w12083 , w12082 , w11119 );
and ( w12084 , w12083 , w11126 );
not ( w12085 , w272 );
and ( w12086 , w12084 , w12085 );
nor ( w12087 , w12086 , w31 );
nor ( w12088 , w12087 , w35 );
nor ( w12089 , w12088 , w37 );
not ( w12090 , w12089 );
and ( w12091 , w12090 , w312 );
not ( w12092 , w12091 );
and ( w12093 , w12092 , w11923 );
nor ( w12094 , w12093 , w12047 );
not ( w12095 , w12063 );
and ( w12096 , w12094 , w12095 );
and ( w12097 , w12096 , w12919 );
not ( w12098 , w12097 );
and ( w12099 , w12098 , w11613 );
not ( w12100 , w12099 );
and ( w12101 , w12100 , g10 );
and ( w12102 , w12101 , g11 );
not ( w12103 , w12102 );
and ( w12104 , w12103 , w11935 );
not ( w12105 , w12104 );
and ( w12106 , w12105 , w11156 );
nor ( w12107 , w12106 , w11094 );
nor ( w12108 , w12107 , w11099 );
nor ( w12109 , w12108 , w11161 );
and ( w12110 , w12109 , w12930 );
nor ( w12111 , w12110 , w53 );
not ( w12112 , w12111 );
and ( w12113 , w12112 , w11285 );
not ( w12114 , w12056 );
and ( w12115 , w12114 , w12113 );
nor ( w12116 , w12115 , w39 );
not ( w12117 , w45 );
and ( w12118 , w12116 , w12117 );
not ( w12119 , w11143 );
and ( w12120 , w12118 , w12119 );
and ( w12121 , w12120 , w11366 );
and ( w12122 , w12121 , w11152 );
and ( w12123 , w12122 , w12919 );
not ( w12124 , w12123 );
and ( w12125 , w12124 , w11613 );
not ( w12126 , w12125 );
and ( w12127 , w12126 , g10 );
and ( w12128 , w12127 , g11 );
not ( w12129 , w12128 );
and ( w12130 , w12129 , w11935 );
not ( w12131 , w12130 );
and ( w12132 , w12131 , w11156 );
nor ( w12133 , w12132 , w11094 );
nor ( w12134 , w12133 , w11099 );
nor ( w12135 , w12134 , w11161 );
and ( w12136 , w12135 , w12930 );
nor ( w12137 , w12136 , w53 );
not ( w12138 , w12137 );
and ( w12139 , w12138 , w11285 );
not ( w12140 , w12048 );
and ( w12141 , w12140 , w12139 );
not ( w12142 , w48 );
and ( w12143 , w12141 , w12142 );
not ( w12144 , w43 );
and ( w12145 , w12143 , w12144 );
nor ( w12146 , w12052 , w12047 );
and ( w12147 , w12146 , w12919 );
not ( w12148 , w12147 );
and ( w12149 , w12148 , w11613 );
not ( w12150 , w12149 );
and ( w12151 , w12150 , g10 );
and ( w12152 , w12151 , g11 );
not ( w12153 , w12152 );
and ( w12154 , w12153 , w11935 );
not ( w12155 , w12154 );
and ( w12156 , w12155 , w11156 );
nor ( w12157 , w12156 , w11094 );
nor ( w12158 , w12157 , w11099 );
nor ( w12159 , w12158 , w11161 );
and ( w12160 , w12159 , w12930 );
nor ( w12161 , w12160 , w53 );
not ( w12162 , w12161 );
and ( w12163 , w12162 , w11285 );
nor ( w12164 , w12145 , w12163 );
and ( w12165 , w12164 , w12919 );
not ( w12166 , w12165 );
and ( w12167 , w12166 , w11613 );
and ( w12168 , w12167 , w11935 );
not ( w12169 , w12168 );
and ( w12170 , w12169 , w11156 );
nor ( w12171 , w12170 , w11094 );
nor ( w12172 , w12171 , w11099 );
nor ( w12173 , w12172 , w11161 );
and ( w12174 , w12173 , w12930 );
nor ( w12175 , w12174 , w53 );
not ( w12176 , w12175 );
and ( w12177 , w12176 , w11285 );
nor ( w12178 , w12047 , w12177 );
and ( w12179 , w12178 , w12560 );
nor ( w12180 , w12063 , w11923 );
nor ( w12181 , w12179 , w12180 );
and ( w12182 , w12181 , w11903 );
not ( w12183 , w12182 );
and ( w12184 , w12183 , g10 );
and ( w12185 , w12184 , g11 );
not ( w12186 , w12185 );
and ( w12187 , w12186 , w11935 );
and ( w12188 , w12187 , w12947 );
nor ( w12189 , w12188 , w53 );
not ( w12190 , w12189 );
and ( w12191 , w12190 , w11285 );
nor ( w12192 , w310 , w12191 );
and ( w12193 , w12192 , w48 );
nor ( w12194 , w12030 , w12191 );
not ( w12195 , w11119 );
and ( w12196 , w12194 , w12195 );
and ( w12197 , w12196 , g30 );
and ( w12198 , w12196 , w12717 );
not ( w12199 , g30 );
and ( w12200 , w12198 , w12199 );
and ( w12201 , w12200 , w12921 );
not ( w12202 , w12201 );
and ( w12203 , w12202 , w11626 );
not ( w12204 , w12203 );
and ( w12205 , w12204 , w11156 );
nor ( w12206 , w12205 , w11094 );
nor ( w12207 , w12206 , w11099 );
nor ( w12208 , w12207 , w11161 );
and ( w12209 , w12208 , w12930 );
nor ( w12210 , w12209 , w53 );
not ( w12211 , w12210 );
and ( w12212 , w12211 , w11285 );
not ( w12213 , w12197 );
and ( w12214 , w12213 , w12212 );
nor ( w12215 , w12214 , w20 );
not ( w12216 , w12215 );
and ( w12217 , w12216 , w11626 );
not ( w12218 , w12217 );
and ( w12219 , w12218 , w11156 );
nor ( w12220 , w12219 , w11094 );
nor ( w12221 , w12220 , w11099 );
nor ( w12222 , w12221 , w11161 );
and ( w12223 , w12222 , w12930 );
nor ( w12224 , w12223 , w53 );
not ( w12225 , w12224 );
and ( w12226 , w12225 , w11285 );
nor ( w12227 , w310 , w12226 );
not ( w12228 , w12227 );
and ( w12229 , w12228 , w12212 );
nor ( w12230 , w12229 , w12051 );
and ( w12231 , w12180 , w377 );
and ( w12232 , w11613 , g10 );
and ( w12233 , w12232 , g11 );
nor ( w12234 , w12233 , w11287 );
and ( w12235 , w12725 , w11819 );
and ( w12236 , w12235 , w12950 );
nor ( w12237 , w12236 , w11099 );
nor ( w12238 , w11104 , w11273 );
and ( w12239 , w12238 , w12950 );
nor ( w12240 , w12239 , w11099 );
and ( w12241 , w12240 , w12612 );
nor ( w12242 , w12237 , w12241 );
and ( w12243 , w12242 , w12930 );
nor ( w12244 , w12243 , w53 );
not ( w12245 , w12244 );
and ( w12246 , w12245 , w11285 );
not ( w12247 , w12234 );
and ( w12248 , w12247 , w12246 );
and ( w12249 , w12248 , w12950 );
nor ( w12250 , w12249 , w11099 );
nor ( w12251 , w12250 , w12241 );
and ( w12252 , w12251 , w12930 );
nor ( w12253 , w12252 , w53 );
not ( w12254 , w12253 );
and ( w12255 , w12254 , w11285 );
nor ( w12256 , w12255 , w11637 );
nor ( w12257 , w12256 , w11094 );
nor ( w12258 , w12257 , w11099 );
and ( w12259 , w12258 , w12612 );
not ( w12260 , w12259 );
and ( w12261 , w12260 , w11285 );
and ( w12262 , w12261 , w12950 );
nor ( w12263 , w12262 , w11099 );
and ( w12264 , w12263 , w12612 );
not ( w12265 , w12264 );
and ( w12266 , w12265 , w11285 );
nor ( w12267 , w12266 , w11637 );
nor ( w12268 , w11114 , w11119 );
and ( w12269 , w12268 , w377 );
nor ( w12270 , w12269 , w11149 );
nor ( w12271 , w11114 , w11119 );
and ( w12272 , w12271 , w377 );
nor ( w12273 , w12272 , w11149 );
and ( w12274 , w12273 , w11670 );
not ( w12275 , w12274 );
and ( w12276 , w12275 , w11174 );
nor ( w12277 , w12276 , w11149 );
not ( w12278 , w12277 );
and ( w12279 , w12278 , w11156 );
nor ( w12280 , w12279 , w11094 );
nor ( w12281 , w12280 , w11099 );
nor ( w12282 , w12281 , w11273 );
nor ( w12283 , w12282 , w53 );
not ( w12284 , w12283 );
and ( w12285 , w12270 , w12284 );
not ( w12286 , w12285 );
and ( w12287 , w12286 , w11174 );
nor ( w12288 , w12287 , w11149 );
not ( w12289 , w12288 );
and ( w12290 , w12289 , w11156 );
nor ( w12291 , w12290 , w11094 );
nor ( w12292 , w12291 , w11099 );
nor ( w12293 , w12292 , w11273 );
nor ( w12294 , w12293 , w53 );
nor ( w12295 , w12294 , w11300 );
not ( w12296 , w12295 );
and ( w12297 , w12296 , w11361 );
and ( w12298 , w12297 , w11366 );
not ( w12299 , w12298 );
and ( w12300 , w12299 , w11285 );
and ( w12301 , w12300 , w12725 );
nor ( w12302 , w12301 , w20 );
nor ( w12303 , w12302 , w11094 );
nor ( w12304 , w12303 , w11099 );
nor ( w12305 , w12304 , w11161 );
and ( w12306 , w12305 , w12905 );
and ( w12307 , w12306 , w12930 );
nor ( w12308 , w12307 , w53 );
not ( w12309 , w12308 );
and ( w12310 , w12309 , w11285 );
and ( w12311 , w12310 , w12905 );
and ( w12312 , w12311 , w11285 );
not ( w12313 , w12267 );
and ( w12314 , w12313 , w12312 );
and ( w12315 , w12314 , w12950 );
and ( w12316 , w12315 , w11285 );
nor ( w12317 , w12316 , w11099 );
and ( w12318 , w12717 , w377 );
and ( w12319 , w12720 , w377 );
nor ( w12320 , w12319 , w11149 );
and ( w12321 , w12320 , w11670 );
and ( w12322 , w12321 , w12725 );
nor ( w12323 , w12322 , w48 );
and ( w12324 , w11285 , w11292 );
and ( w12325 , w12324 , w12725 );
and ( w12326 , w12325 , w11285 );
and ( w12327 , w12326 , w11630 );
and ( w12328 , w12327 , w11285 );
and ( w12329 , w12328 , w11630 );
and ( w12330 , w11285 , w12329 );
nor ( w12331 , w11291 , w11300 );
and ( w12332 , w12331 , w12725 );
and ( w12333 , w12330 , w12332 );
and ( w12334 , w12333 , w12725 );
and ( w12335 , w12334 , w11285 );
and ( w12336 , w12335 , w12725 );
and ( w12337 , w12336 , w12950 );
nor ( w12338 , w12337 , w11099 );
nor ( w12339 , w12338 , w11161 );
and ( w12340 , w12339 , w12905 );
and ( w12341 , w12340 , w12930 );
nor ( w12342 , w12341 , w53 );
not ( w12343 , w12342 );
and ( w12344 , w12343 , w11285 );
not ( w12345 , w12323 );
and ( w12346 , w12345 , w12344 );
not ( w12347 , w12346 );
and ( w12348 , w12347 , w11275 );
and ( w12349 , w12348 , w11156 );
nor ( w12350 , w12349 , w11094 );
nor ( w12351 , w12350 , w11099 );
nor ( w12352 , w12351 , w11161 );
and ( w12353 , w12352 , w12905 );
and ( w12354 , w12353 , w12930 );
nor ( w12355 , w12354 , w53 );
not ( w12356 , w12355 );
and ( w12357 , w12356 , w11285 );
not ( w12358 , w12318 );
and ( w12359 , w12358 , w12357 );
nor ( w12360 , w12359 , w12051 );
and ( w12361 , w12344 , w11670 );
nor ( w12362 , w11903 , w11114 );
not ( w12363 , w12362 );
and ( w12364 , w12363 , w11630 );
and ( w12365 , w12364 , w11670 );
and ( w12366 , w12365 , w12725 );
and ( w12367 , w12366 , w12344 );
and ( w12368 , w12367 , w12950 );
nor ( w12369 , w12368 , w11099 );
nor ( w12370 , w12369 , w11161 );
and ( w12371 , w12370 , w12905 );
nor ( w12372 , w12371 , w53 );
not ( w12373 , w12372 );
and ( w12374 , w12373 , w11285 );
and ( w12375 , w12255 , w12374 );
nor ( w12376 , w624 , w11099 );
and ( w12377 , w12376 , w12612 );
and ( w12378 , w12375 , w12764 );
not ( w12379 , g34 );
and ( w12380 , w12378 , w12379 );
not ( w12381 , g35 );
and ( w12382 , w12380 , w12381 );
and ( w12383 , w12329 , w12332 );
and ( w12384 , w12383 , w11285 );
and ( w12385 , w12384 , w12725 );
and ( w12386 , w12385 , w11285 );
and ( w12387 , w12386 , w12725 );
and ( w12388 , w12387 , w7791 );
and ( w12389 , w7791 , w13211 );
nor ( w12390 , w12389 , w53 );
not ( w12391 , w12390 );
and ( w12392 , w12391 , w11285 );
and ( w12393 , w7791 , w12392 );
and ( w12394 , w12393 , w12725 );
and ( w12395 , w12394 , w11630 );
and ( w12396 , w12395 , w12950 );
nor ( w12397 , w12396 , w11099 );
and ( w12398 , w12397 , w12612 );
not ( w12399 , w12398 );
and ( w12400 , w12399 , w11285 );
and ( w12401 , w12388 , w12400 );
and ( w12402 , w12401 , w12725 );
and ( w12403 , w12402 , w11630 );
and ( w12404 , w12403 , w12950 );
nor ( w12405 , w12404 , w11099 );
nor ( w12406 , w12405 , w11161 );
and ( w12407 , w12406 , w12905 );
and ( w12408 , w12407 , w12930 );
nor ( w12409 , w12408 , w53 );
not ( w12410 , w12409 );
and ( w12411 , w12410 , w11285 );
not ( w12412 , w12411 );
and ( w12413 , w12412 , w308 );
nor ( w12414 , g35 , w349 );
nor ( w12415 , w12413 , w12414 );
and ( w12416 , w12415 , w12266 );
and ( w12417 , w12416 , w12344 );
and ( w12418 , w12417 , w11670 );
and ( w12419 , w12418 , w11630 );
and ( w12420 , w12419 , w11626 );
and ( w12421 , w12420 , w12725 );
nor ( w12422 , w12421 , w11637 );
and ( w12423 , w11831 , w12725 );
not ( w12424 , w37 );
and ( w12425 , w12328 , w12424 );
and ( w12426 , w12425 , w11630 );
nor ( w12427 , w12426 , w39 );
not ( w12428 , w12427 );
and ( w12429 , w12428 , w11285 );
nor ( w12430 , w12429 , w45 );
not ( w12431 , w12430 );
and ( w12432 , w12431 , w11285 );
and ( w12433 , w12432 , w12332 );
and ( w12434 , w12433 , w12725 );
nor ( w12435 , w12434 , w11099 );
nor ( w12436 , w12435 , w11161 );
nor ( w12437 , w12436 , w53 );
not ( w12438 , w12437 );
and ( w12439 , w12438 , w11285 );
and ( w12440 , w11670 , w12439 );
and ( w12441 , w12440 , w11285 );
nor ( w12442 , w12441 , w18 );
nor ( w12443 , w12442 , w11149 );
and ( w12444 , w20 , w12612 );
not ( w12445 , w12444 );
and ( w12446 , w12443 , w12445 );
nor ( w12447 , w12446 , w11287 );
not ( w12448 , w12447 );
and ( w12449 , w12448 , w11831 );
and ( w12450 , w12449 , w12725 );
and ( w12451 , w12446 , w12725 );
nor ( w12452 , w12451 , w11287 );
not ( w12453 , w12452 );
and ( w12454 , w12453 , w11831 );
and ( w12455 , w12454 , w12950 );
nor ( w12456 , w12455 , w11099 );
nor ( w12457 , w12456 , w11161 );
and ( w12458 , w12457 , w12930 );
nor ( w12459 , w12458 , w53 );
not ( w12460 , w12459 );
and ( w12461 , w12460 , w11285 );
and ( w12462 , w12450 , w12461 );
and ( w12463 , w12462 , w12725 );
nor ( w12464 , w12463 , w19 );
and ( w12465 , w12464 , w11156 );
nor ( w12466 , w12465 , w11094 );
nor ( w12467 , w12466 , w11099 );
nor ( w12468 , w12467 , w11161 );
and ( w12469 , w12468 , w12905 );
and ( w12470 , w12469 , w12930 );
nor ( w12471 , w12470 , w53 );
not ( w12472 , w12471 );
and ( w12473 , w12472 , w11285 );
and ( w12474 , w12423 , w12473 );
and ( w12475 , w12474 , w12947 );
and ( w12476 , w12475 , w11285 );
not ( w12477 , w12422 );
and ( w12478 , w12477 , w12476 );
and ( w12479 , w12478 , w12950 );
nor ( w12480 , w12479 , w11099 );
nor ( w12481 , w12480 , w11273 );
nor ( w12482 , w12481 , w53 );
not ( w12483 , w12482 );
and ( w12484 , w12483 , w11285 );
and ( w12485 , w12361 , w12484 );
and ( w12486 , w12485 , w11630 );
and ( w12487 , w12486 , w11626 );
and ( w12488 , w12487 , w12725 );
nor ( w12489 , w12488 , w11637 );
not ( w12490 , w12489 );
and ( w12491 , w12490 , w12476 );
and ( w12492 , w12491 , w12950 );
nor ( w12493 , w12492 , w11099 );
nor ( w12494 , w12493 , w11273 );
nor ( w12495 , w12494 , w53 );
not ( w12496 , w12495 );
and ( w12497 , w12496 , w11285 );
not ( w12498 , w377 );
and ( w12499 , w12498 , w12497 );
and ( w12500 , w12344 , w11114 );
and ( w12501 , w12500 , g30 );
and ( w12502 , w12501 , g31 );
not ( w12503 , w12502 );
and ( w12504 , w12503 , w377 );
not ( w12505 , w12504 );
and ( w12506 , w12505 , w12497 );
and ( w12507 , w12506 , w11626 );
nor ( w12508 , w12507 , w11637 );
not ( w12509 , w12508 );
and ( w12510 , w12509 , w12476 );
and ( w12511 , w12510 , w12950 );
nor ( w12512 , w12511 , w11099 );
nor ( w12513 , w12512 , w11273 );
nor ( w12514 , w12513 , w53 );
not ( w12515 , w12514 );
and ( w12516 , w12515 , w11285 );
not ( w12517 , w12516 );
and ( w12518 , w12517 , w308 );
not ( w12519 , w12518 );
and ( w12520 , w12519 , w12392 );
not ( w12521 , w12520 );
and ( w12522 , w12521 , w308 );
and ( w12523 , w12231 , w13536 );
and ( w12524 , w12523 , w12612 );
not ( w12525 , w12524 );
and ( w12526 , w12525 , w11285 );
not ( w12527 , w12414 );
and ( w12528 , w12526 , w12527 );
not ( w12529 , w11109 );
and ( w12530 , g30 , w12529 );
nor ( w12531 , w12530 , w12051 );
not ( w12532 , w308 );
and ( w12533 , w12052 , w12532 );
nor ( w12534 , w12533 , w53 );
not ( w12535 , w12534 );
and ( w12536 , w12535 , w11285 );
nor ( w12537 , w12536 , g30 );
nor ( w12538 , w12537 , w11109 );
not ( w12539 , w12536 );
and ( w12540 , w12539 , w11156 );
nor ( w12541 , w12540 , w11094 );
nor ( w12542 , w12541 , w11099 );
nor ( w12543 , w12542 , w11273 );
nor ( w12544 , w12543 , w53 );
not ( w12545 , w12544 );
and ( w12546 , w12545 , w11285 );
nor ( w12547 , w12538 , w12546 );
nor ( w12548 , w12547 , w12180 );
nor ( w12549 , w12548 , w7791 );
and ( w12550 , w12549 , w11156 );
nor ( w12551 , w12550 , w11094 );
nor ( w12552 , w12551 , w11099 );
nor ( w12553 , w12552 , w11273 );
nor ( w12554 , w12553 , w53 );
not ( w12555 , w12554 );
and ( w12556 , w12555 , w11285 );
not ( w12557 , w12531 );
and ( w12558 , w12557 , w12556 );
nor ( w12559 , w11114 , w12139 );
not ( w12560 , w12051 );
and ( w12561 , w12559 , w12560 );
not ( w12562 , w7791 );
and ( w12563 , w12559 , w12562 );
not ( w12564 , w12563 );
and ( w12565 , w12564 , w11847 );
and ( w12566 , w12565 , w12725 );
not ( w12567 , w12566 );
and ( w12568 , w12567 , w11156 );
nor ( w12569 , w12568 , w11094 );
nor ( w12570 , w12569 , w11099 );
nor ( w12571 , w12570 , w11273 );
nor ( w12572 , w12571 , w53 );
not ( w12573 , w12572 );
and ( w12574 , w12573 , w11285 );
not ( w12575 , w12561 );
and ( w12576 , w12575 , w12574 );
and ( w12577 , w12576 , w11285 );
and ( w12578 , w12577 , w12725 );
and ( w12579 , w12578 , w12344 );
not ( w12580 , w12579 );
and ( w12581 , w12580 , w11275 );
nor ( w12582 , w12581 , w11149 );
and ( w12583 , w12582 , w12950 );
nor ( w12584 , w12583 , w11099 );
nor ( w12585 , w12584 , w11161 );
and ( w12586 , w12585 , w12905 );
and ( w12587 , w12586 , w12930 );
nor ( w12588 , w12587 , w53 );
not ( w12589 , w12588 );
and ( w12590 , w12589 , w11285 );
and ( w12591 , w12558 , w12590 );
not ( w12592 , w12591 );
and ( w12593 , w12592 , w377 );
not ( w12594 , w12593 );
and ( w12595 , w12594 , w12497 );
not ( w12596 , w12595 );
and ( w12597 , w12596 , w11275 );
not ( w12598 , w12597 );
and ( w12599 , w12598 , w11626 );
and ( w12600 , w12599 , w12725 );
nor ( w12601 , w12600 , w11637 );
not ( w12602 , w12601 );
and ( w12603 , w12602 , w12476 );
and ( w12604 , w12603 , w12950 );
nor ( w12605 , w12604 , w11099 );
nor ( w12606 , w12605 , w11273 );
nor ( w12607 , w12606 , w53 );
not ( w12608 , w12607 );
and ( w12609 , w12608 , w11285 );
and ( w12610 , w12609 , w12950 );
nor ( w12611 , w12610 , w11099 );
not ( w12612 , w53 );
and ( w12613 , w12611 , w12612 );
not ( w12614 , w12613 );
and ( w12615 , w12614 , w11285 );
and ( w12616 , w12344 , w12615 );
and ( w12617 , w12616 , w12497 );
and ( w12618 , w12617 , w11626 );
nor ( w12619 , w12618 , w11637 );
not ( w12620 , w12619 );
and ( w12621 , w12620 , w12476 );
and ( w12622 , w12621 , w12950 );
nor ( w12623 , w12622 , w11099 );
nor ( w12624 , w12623 , w11273 );
nor ( w12625 , w12624 , w53 );
not ( w12626 , w12625 );
and ( w12627 , w12626 , w11285 );
and ( w12628 , w12528 , w12627 );
nor ( w12629 , w12628 , w53 );
not ( w12630 , w12629 );
and ( w12631 , w12630 , w11285 );
not ( w12632 , w12522 );
and ( w12633 , w12632 , w12631 );
not ( w12634 , w12633 );
and ( w12635 , w12634 , w11275 );
not ( w12636 , w12635 );
and ( w12637 , w12636 , w11626 );
nor ( w12638 , w12637 , w11637 );
not ( w12639 , w12638 );
and ( w12640 , w12639 , w12476 );
and ( w12641 , w12640 , w12950 );
nor ( w12642 , w12641 , w11099 );
nor ( w12643 , w12642 , w11273 );
nor ( w12644 , w12643 , w53 );
not ( w12645 , w12644 );
and ( w12646 , w12645 , w11285 );
nor ( w12647 , w12499 , w12646 );
and ( w12648 , w12647 , w11275 );
not ( w12649 , w12648 );
and ( w12650 , w12649 , w11626 );
nor ( w12651 , w12650 , w11637 );
not ( w12652 , w11305 );
and ( w12653 , w12652 , w12344 );
and ( w12654 , w12653 , w12725 );
and ( w12655 , w12654 , w12950 );
nor ( w12656 , w12655 , w11099 );
nor ( w12657 , w12656 , w11161 );
and ( w12658 , w12657 , w12905 );
and ( w12659 , w12658 , w12930 );
nor ( w12660 , w12659 , w53 );
not ( w12661 , w12660 );
and ( w12662 , w12661 , w11285 );
and ( w12663 , w11670 , w12662 );
and ( w12664 , w12663 , w11285 );
and ( w12665 , w12664 , w12725 );
and ( w12666 , w12665 , w12950 );
nor ( w12667 , w12666 , w11099 );
nor ( w12668 , w12667 , w11273 );
nor ( w12669 , w12668 , w53 );
not ( w12670 , w12669 );
and ( w12671 , w12670 , w11285 );
and ( w12672 , w12671 , w11630 );
and ( w12673 , w12672 , w12725 );
and ( w12674 , w12673 , w11831 );
and ( w12675 , w12674 , w12947 );
and ( w12676 , w12675 , w12905 );
and ( w12677 , w12676 , w11285 );
not ( w12678 , w12651 );
and ( w12679 , w12678 , w12677 );
and ( w12680 , w12679 , w12950 );
nor ( w12681 , w12680 , w11099 );
nor ( w12682 , w12681 , w11273 );
nor ( w12683 , w12682 , w53 );
not ( w12684 , w12683 );
and ( w12685 , w12684 , w11285 );
nor ( w12686 , w12382 , w12685 );
not ( w12687 , w12686 );
and ( w12688 , w12687 , w11626 );
and ( w12689 , w12688 , w11630 );
nor ( w12690 , w12689 , w11637 );
not ( w12691 , w12690 );
and ( w12692 , w12691 , w12677 );
and ( w12693 , w12692 , w12950 );
nor ( w12694 , w12693 , w11099 );
nor ( w12695 , w12694 , w11273 );
nor ( w12696 , w12695 , w53 );
not ( w12697 , w12696 );
and ( w12698 , w12697 , w11285 );
and ( w12699 , w12361 , w12698 );
and ( w12700 , w12699 , w11847 );
and ( w12701 , w12700 , w12764 );
nor ( w12702 , w12701 , w12685 );
not ( w12703 , w12702 );
and ( w12704 , w12703 , w11626 );
and ( w12705 , w12704 , w11630 );
nor ( w12706 , w12705 , w11637 );
not ( w12707 , w12706 );
and ( w12708 , w12707 , w12677 );
and ( w12709 , w12708 , w12950 );
nor ( w12710 , w12709 , w11099 );
nor ( w12711 , w12710 , w11273 );
nor ( w12712 , w12711 , w53 );
not ( w12713 , w12712 );
and ( w12714 , w12713 , w11285 );
not ( w12715 , w12360 );
and ( w12716 , w12715 , w12714 );
not ( w12717 , w310 );
and ( w12718 , w12717 , w308 );
and ( w12719 , w12718 , w377 );
not ( w12720 , w11114 );
and ( w12721 , w308 , w12720 );
and ( w12722 , w12721 , w377 );
nor ( w12723 , w12722 , w11149 );
and ( w12724 , w12723 , w11670 );
not ( w12725 , w11149 );
and ( w12726 , w12724 , w12725 );
nor ( w12727 , w12726 , w48 );
not ( w12728 , w12727 );
and ( w12729 , w12728 , w12344 );
not ( w12730 , w12729 );
and ( w12731 , w12730 , w308 );
and ( w12732 , w12731 , w11275 );
and ( w12733 , w12732 , w11156 );
nor ( w12734 , w12733 , w11094 );
nor ( w12735 , w12734 , w11099 );
nor ( w12736 , w12735 , w11161 );
and ( w12737 , w12736 , w12905 );
and ( w12738 , w12737 , w12930 );
nor ( w12739 , w12738 , w53 );
not ( w12740 , w12739 );
and ( w12741 , w12740 , w11285 );
not ( w12742 , w12719 );
and ( w12743 , w12742 , w12741 );
not ( w12744 , w12743 );
and ( w12745 , w12744 , w308 );
nor ( w12746 , w12745 , w12377 );
nor ( w12747 , w12746 , w12685 );
and ( w12748 , w12747 , w11275 );
and ( w12749 , w12748 , w12919 );
not ( w12750 , w12749 );
and ( w12751 , w12750 , w11626 );
and ( w12752 , w12751 , w11630 );
nor ( w12753 , w12752 , w11637 );
not ( w12754 , w12753 );
and ( w12755 , w12754 , w12677 );
and ( w12756 , w12755 , w12950 );
nor ( w12757 , w12756 , w11099 );
nor ( w12758 , w12757 , w11161 );
and ( w12759 , w12758 , w12930 );
nor ( w12760 , w12759 , w53 );
not ( w12761 , w12760 );
and ( w12762 , w12761 , w11285 );
and ( w12763 , w12716 , w12762 );
not ( w12764 , w12377 );
and ( w12765 , w12763 , w12764 );
nor ( w12766 , w12765 , w12685 );
and ( w12767 , w12766 , w11275 );
and ( w12768 , w12767 , w12919 );
not ( w12769 , w12768 );
and ( w12770 , w12769 , w11626 );
and ( w12771 , w12770 , w11630 );
nor ( w12772 , w12771 , w11637 );
not ( w12773 , w12772 );
and ( w12774 , w12773 , w12677 );
and ( w12775 , w12774 , w12950 );
nor ( w12776 , w12775 , w11099 );
nor ( w12777 , w12776 , w11161 );
and ( w12778 , w12777 , w12930 );
nor ( w12779 , w12778 , w53 );
not ( w12780 , w12779 );
and ( w12781 , w12780 , w11285 );
not ( w12782 , w12317 );
and ( w12783 , w12782 , w12781 );
and ( w12784 , w12783 , w12905 );
nor ( w12785 , w12784 , w53 );
not ( w12786 , w12785 );
and ( w12787 , w12786 , w11630 );
not ( w12788 , w12392 );
and ( w12789 , w12788 , w308 );
not ( w12790 , w12789 );
and ( w12791 , w12790 , w12526 );
nor ( w12792 , w12791 , w53 );
not ( w12793 , w12792 );
and ( w12794 , w12793 , w11285 );
and ( w12795 , w12787 , w12794 );
and ( w12796 , w12795 , w11285 );
not ( w12797 , w12231 );
and ( w12798 , w12797 , w12796 );
and ( w12799 , w12798 , w12312 );
and ( w12800 , w12799 , w12950 );
and ( w12801 , w12800 , w11285 );
nor ( w12802 , w12801 , w11099 );
not ( w12803 , w12802 );
and ( w12804 , w12803 , w12781 );
and ( w12805 , w12804 , w12905 );
nor ( w12806 , w12805 , w53 );
not ( w12807 , w12806 );
and ( w12808 , w12807 , w11630 );
and ( w12809 , w12808 , w12794 );
and ( w12810 , w12809 , w11285 );
not ( w12811 , w12230 );
and ( w12812 , w12811 , w12810 );
not ( w12813 , w12812 );
and ( w12814 , w12813 , w377 );
not ( w12815 , w12814 );
and ( w12816 , w12815 , w12796 );
nor ( w12817 , w12816 , w18 );
not ( w12818 , w12817 );
and ( w12819 , w12818 , w11626 );
nor ( w12820 , w12819 , w11637 );
not ( w12821 , w12820 );
and ( w12822 , w12821 , w12312 );
not ( w12823 , w12822 );
and ( w12824 , w12823 , w11174 );
nor ( w12825 , w12824 , w11094 );
and ( w12826 , w12825 , w11285 );
not ( w12827 , w12826 );
and ( w12828 , w12827 , w41 );
and ( w12829 , w12828 , w13536 );
not ( w12830 , w12829 );
and ( w12831 , w12830 , w12781 );
and ( w12832 , w12831 , w12947 );
and ( w12833 , w12832 , w12905 );
and ( w12834 , w12833 , w12930 );
nor ( w12835 , w12834 , w53 );
not ( w12836 , w12835 );
and ( w12837 , w12836 , w11630 );
and ( w12838 , w12837 , w12794 );
and ( w12839 , w12838 , w11285 );
not ( w12840 , w12193 );
and ( w12841 , w12840 , w12839 );
nor ( w12842 , w12841 , w12051 );
not ( w12843 , w12842 );
and ( w12844 , w12843 , w12810 );
not ( w12845 , w12844 );
and ( w12846 , w12845 , w377 );
not ( w12847 , w12846 );
and ( w12848 , w12847 , w12796 );
nor ( w12849 , w12848 , w11637 );
not ( w12850 , w12849 );
and ( w12851 , w12850 , w12312 );
not ( w12852 , w12851 );
and ( w12853 , w12852 , w11156 );
nor ( w12854 , w12853 , w11094 );
and ( w12855 , w12854 , w11285 );
not ( w12856 , w12855 );
and ( w12857 , w12856 , w41 );
and ( w12858 , w12857 , w13536 );
not ( w12859 , w12858 );
and ( w12860 , w12859 , w12781 );
and ( w12861 , w12860 , w12905 );
and ( w12862 , w12861 , w12930 );
nor ( w12863 , w12862 , w53 );
not ( w12864 , w12863 );
and ( w12865 , w12864 , w11630 );
and ( w12866 , w12865 , w12794 );
and ( w12867 , w12866 , w11285 );
not ( w12868 , w12036 );
and ( w12869 , w12868 , w12867 );
not ( w12870 , w12869 );
and ( w12871 , w12870 , w377 );
not ( w12872 , w12871 );
and ( w12873 , w12872 , w12796 );
nor ( w12874 , w12873 , w18 );
and ( w12875 , w12874 , w12921 );
not ( w12876 , w12875 );
and ( w12877 , w12876 , w11626 );
nor ( w12878 , w12877 , w11637 );
not ( w12879 , w12878 );
and ( w12880 , w12879 , w12312 );
not ( w12881 , w12880 );
and ( w12882 , w12881 , w11156 );
and ( w12883 , w12882 , w11174 );
nor ( w12884 , w12883 , w11094 );
and ( w12885 , w12884 , w11285 );
not ( w12886 , w12885 );
and ( w12887 , w12886 , w41 );
and ( w12888 , w12887 , w13536 );
not ( w12889 , w12888 );
and ( w12890 , w12889 , w12781 );
and ( w12891 , w12890 , w12947 );
and ( w12892 , w12891 , w12905 );
and ( w12893 , w12892 , w12930 );
nor ( w12894 , w12893 , w53 );
not ( w12895 , w12894 );
and ( w12896 , w12895 , w11630 );
and ( w12897 , w12896 , w12794 );
and ( w12898 , w12897 , w11285 );
and ( w12899 , w12898 , w12312 );
and ( w12900 , w12899 , w12950 );
and ( w12901 , w12900 , w11285 );
nor ( w12902 , w12901 , w11099 );
not ( w12903 , w12902 );
and ( w12904 , w12903 , w12781 );
not ( w12905 , w12241 );
and ( w12906 , w12904 , w12905 );
nor ( w12907 , w12906 , w53 );
not ( w12908 , w12907 );
and ( w12909 , w12908 , w11630 );
and ( w12910 , w12909 , w12794 );
and ( w12911 , w12910 , w11285 );
not ( w12912 , w12029 );
and ( w12913 , w12912 , w12911 );
and ( w12914 , w12913 , w12950 );
and ( w12915 , w12914 , w12018 );
nor ( w12916 , w12915 , w11099 );
nor ( w12917 , w12916 , w11104 );
nor ( w12918 , w12917 , w53 );
not ( w12919 , w18 );
and ( w12920 , w12918 , w12919 );
not ( w12921 , w20 );
and ( w12922 , w12920 , w12921 );
not ( w12923 , w12922 );
and ( w12924 , w12923 , w11626 );
nor ( w12925 , w12924 , w11637 );
nor ( w12926 , w12925 , w11094 );
and ( w12927 , w12926 , w12018 );
nor ( w12928 , w12927 , w11099 );
nor ( w12929 , w12928 , w11104 );
not ( w12930 , w11273 );
and ( w12931 , w12929 , w12930 );
nor ( w12932 , w12931 , w53 );
nor ( w12933 , w224 , w218 );
not ( w12934 , g7 );
and ( w12935 , w12933 , w12934 );
and ( w12936 , w12935 , w13536 );
and ( w12937 , w12936 , w11094 );
nor ( w12938 , w12937 , w11284 );
not ( w12939 , w12932 );
and ( w12940 , w12939 , w12938 );
and ( w12941 , w12940 , w12911 );
and ( w12942 , w12941 , w12018 );
and ( w12943 , w12942 , w13367 );
and ( w12944 , w12943 , w12938 );
and ( w12945 , w12944 , g48 );
and ( w12946 , w12945 , g31 );
not ( w12947 , w11161 );
and ( w12948 , w12947 , w12944 );
and ( w12949 , w13584 , w12948 );
not ( w12950 , w11094 );
and ( w12951 , w12950 , w12949 );
nor ( w12952 , w11099 , w12951 );
not ( w12953 , w12946 );
and ( w12954 , w12953 , w12952 );
and ( w12955 , w13607 , g41 );
and ( w12956 , w12955 , g15 );
and ( w12957 , w12956 , w13607 );
not ( w12958 , w12957 );
and ( w12959 , w12958 , w12948 );
not ( w12960 , w12959 );
and ( w12961 , w12960 , w12952 );
not ( w12962 , g38 );
and ( w12963 , g25 , w12962 );
not ( w12964 , g25 );
and ( w12965 , w12964 , g38 );
and ( w12966 , w12965 , w13536 );
and ( w12967 , w12966 , w11094 );
nor ( w12968 , w12967 , w11284 );
not ( w12969 , w12963 );
and ( w12970 , w12969 , w12968 );
nor ( w12971 , w12970 , g17 );
not ( w12972 , w12971 );
and ( w12973 , w12972 , g40 );
nor ( w12974 , w12970 , w11099 );
and ( w12975 , w12974 , w11094 );
nor ( w12976 , w12975 , w11284 );
nor ( w12977 , w12973 , w12976 );
and ( w12978 , w12977 , w13536 );
and ( w12979 , w12978 , w11094 );
nor ( w12980 , w12979 , w11284 );
not ( w12981 , w12961 );
and ( w12982 , w12981 , w12980 );
and ( w12983 , w12982 , w12948 );
nor ( w12984 , w12983 , w12976 );
not ( w12985 , w12984 );
and ( w12986 , w12985 , w12948 );
and ( w12987 , w12986 , w11718 );
and ( w12988 , w12987 , w12948 );
nor ( w12989 , w12988 , w12951 );
and ( w12990 , w12989 , w12952 );
and ( w12991 , w12990 , g25 );
not ( w12992 , w12968 );
and ( w12993 , w12992 , g38 );
and ( w12994 , w12993 , w13536 );
and ( w12995 , w12994 , w11094 );
nor ( w12996 , w12995 , w11284 );
nor ( w12997 , w12996 , w12968 );
and ( w12998 , w12997 , g38 );
and ( w12999 , w12998 , w13536 );
and ( w13000 , w12999 , w11094 );
nor ( w13001 , w13000 , w11284 );
nor ( w13002 , w13001 , g25 );
and ( w13003 , w13002 , g38 );
and ( w13004 , w13003 , w13536 );
and ( w13005 , w13004 , w11094 );
nor ( w13006 , w13005 , w11284 );
not ( w13007 , w12991 );
and ( w13008 , w13007 , w13006 );
and ( w13009 , w13008 , w12948 );
nor ( w13010 , w13009 , w11722 );
not ( w13011 , w13010 );
and ( w13012 , w13011 , w12948 );
not ( w13013 , w11720 );
and ( w13014 , w13012 , w13013 );
not ( w13015 , w13014 );
and ( w13016 , w13015 , w12952 );
not ( w13017 , w13016 );
and ( w13018 , w13017 , w12944 );
not ( w13019 , w13018 );
and ( w13020 , w13019 , w12952 );
and ( w13021 , w13020 , w13607 );
and ( w13022 , w13021 , w12952 );
and ( w13023 , w12944 , g42 );
and ( w13024 , w13023 , g21 );
nor ( w13025 , w13024 , w12951 );
and ( w13026 , w13022 , w13025 );
and ( w13027 , w13026 , w13536 );
and ( w13028 , w11186 , w13545 );
nor ( w13029 , w13028 , w11099 );
and ( w13030 , w13029 , w11094 );
not ( w13031 , w13030 );
and ( w13032 , w13031 , w12949 );
and ( w13033 , w11817 , w11670 );
and ( w13034 , w13033 , w11819 );
and ( w13035 , w13034 , w13584 );
and ( w13036 , w11819 , w13035 );
and ( w13037 , w13036 , w12948 );
and ( w13038 , w13032 , w13037 );
and ( w13039 , w13038 , w12948 );
not ( w13040 , w13039 );
and ( w13041 , w13027 , w13040 );
not ( w13042 , w11193 );
and ( w13043 , w13042 , w11747 );
nor ( w13044 , w13043 , w11284 );
not ( w13045 , w1934 );
and ( w13046 , w13045 , w11756 );
nor ( w13047 , w13046 , w11193 );
and ( w13048 , w13047 , w11656 );
nor ( w13049 , w11193 , w11756 );
not ( w13050 , g27 );
and ( w13051 , w13050 , g44 );
not ( w13052 , w13051 );
and ( w13053 , w13052 , w11094 );
nor ( w13054 , w13053 , w11284 );
and ( w13055 , w13054 , w13367 );
not ( w13056 , w13055 );
and ( w13057 , g44 , w13056 );
nor ( w13058 , w13057 , w11104 );
nor ( w13059 , w11104 , w11284 );
and ( w13060 , w13058 , w13059 );
and ( w13061 , w13060 , w13367 );
and ( w13062 , w13061 , w13059 );
and ( w13063 , w13062 , w13367 );
and ( w13064 , w13584 , w13063 );
nor ( w13065 , w13064 , w11752 );
nor ( w13066 , w13065 , w11104 );
and ( w13067 , w13066 , w13059 );
not ( w13068 , w13067 );
and ( w13069 , w13068 , w11094 );
nor ( w13070 , w13069 , w11284 );
and ( w13071 , w13070 , w13367 );
not ( w13072 , w13049 );
and ( w13073 , w13072 , w13071 );
and ( w13074 , w13073 , w13584 );
and ( w13075 , w13074 , w11670 );
and ( w13076 , w13075 , w13058 );
and ( w13077 , w13076 , w13367 );
nor ( w13078 , w13077 , w11752 );
nor ( w13079 , w13078 , w11104 );
nor ( w13080 , w13079 , w11758 );
nor ( w13081 , w13080 , w11104 );
nor ( w13082 , w13081 , w11186 );
and ( w13083 , w11670 , w11819 );
and ( w13084 , w13083 , w13584 );
not ( w13085 , w13082 );
and ( w13086 , w13085 , w13084 );
not ( w13087 , w13086 );
and ( w13088 , w13087 , w11094 );
nor ( w13089 , w13088 , w11284 );
and ( w13090 , w13089 , w13367 );
not ( w13091 , w13048 );
and ( w13092 , w13091 , w13090 );
and ( w13093 , w13092 , w13058 );
and ( w13094 , w13093 , w13367 );
nor ( w13095 , w13094 , w11752 );
nor ( w13096 , w13095 , w11104 );
nor ( w13097 , w13096 , w11758 );
nor ( w13098 , w13097 , w11104 );
nor ( w13099 , w13098 , w11186 );
not ( w13100 , w13099 );
and ( w13101 , w13100 , w13084 );
not ( w13102 , w13101 );
and ( w13103 , w13102 , w11094 );
nor ( w13104 , w13103 , w11284 );
and ( w13105 , w13104 , w13367 );
and ( w13106 , w13044 , w13105 );
and ( w13107 , w13106 , w13584 );
and ( w13108 , w13107 , w13367 );
nor ( w13109 , w13108 , g45 );
and ( w13110 , w13109 , w13333 );
and ( w13111 , w13064 , w11670 );
and ( w13112 , w13111 , w13584 );
and ( w13113 , w13112 , w11670 );
nor ( w13114 , w13113 , w11752 );
nor ( w13115 , w13114 , w11104 );
and ( w13116 , w13115 , w13059 );
and ( w13117 , w13116 , w13084 );
not ( w13118 , w13117 );
and ( w13119 , w13118 , w11094 );
nor ( w13120 , w13119 , w11284 );
and ( w13121 , w13120 , w13367 );
not ( w13122 , w13110 );
and ( w13123 , w13122 , w13121 );
and ( w13124 , w13123 , w13367 );
and ( w13125 , w13124 , w13584 );
and ( w13126 , w11783 , w11753 );
and ( w13127 , w13126 , w11199 );
and ( w13128 , w13127 , w11094 );
and ( w13129 , w13125 , w13570 );
nor ( w13130 , w13129 , w11758 );
nor ( w13131 , w13130 , w11104 );
and ( w13132 , w13131 , w13059 );
and ( w13133 , w13084 , w13059 );
and ( w13134 , w13133 , w13367 );
and ( w13135 , w13134 , w13084 );
and ( w13136 , w13135 , w13584 );
and ( w13137 , w13136 , w13367 );
and ( w13138 , w13132 , w13137 );
and ( w13139 , w13138 , w13584 );
nor ( w13140 , w13139 , w11762 );
and ( w13141 , w13140 , w13257 );
nor ( w13142 , w13141 , w11284 );
and ( w13143 , w13142 , w13367 );
and ( w13144 , w13059 , w11817 );
and ( w13145 , w13144 , w13584 );
and ( w13146 , w13145 , w13367 );
and ( w13147 , w13143 , w13146 );
and ( w13148 , w13147 , w13084 );
not ( w13149 , w13148 );
and ( w13150 , w13149 , w11199 );
not ( w13151 , w13150 );
and ( w13152 , w13151 , w13059 );
not ( w13153 , w13152 );
and ( w13154 , w13153 , w11094 );
nor ( w13155 , w13154 , w11284 );
and ( w13156 , w13155 , w13367 );
and ( w13157 , w13156 , w13084 );
and ( w13158 , w13157 , w13367 );
and ( w13159 , w13158 , w12911 );
nor ( w13160 , w9711 , w9108 );
nor ( w13161 , w11728 , w11099 );
and ( w13162 , g41 , g15 );
not ( w13163 , w12976 );
and ( w13164 , w13162 , w13163 );
not ( w13165 , w13164 );
and ( w13166 , w13165 , w12980 );
and ( w13167 , w13166 , w11718 );
and ( w13168 , w13167 , g25 );
nor ( w13169 , w13168 , g38 );
not ( w13170 , w13169 );
and ( w13171 , w13170 , w13006 );
and ( w13172 , w13171 , w13584 );
and ( w13173 , w13172 , w13503 );
nor ( w13174 , w13173 , w11193 );
and ( w13175 , w13059 , w12911 );
not ( w13176 , w13174 );
and ( w13177 , w13176 , w13175 );
nor ( w13178 , w11193 , w11099 );
and ( w13179 , w11653 , w13536 );
and ( w13180 , w13179 , w11094 );
nor ( w13181 , w13180 , w11284 );
and ( w13182 , w13181 , w13367 );
nor ( w13183 , w13182 , g31 );
nor ( w13184 , w13183 , g45 );
and ( w13185 , w13184 , w13333 );
not ( w13186 , w13185 );
and ( w13187 , w13186 , g48 );
nor ( w13188 , w13182 , g29 );
and ( w13189 , w13188 , w13204 );
and ( w13190 , w13189 , w13536 );
and ( w13191 , w13190 , w11094 );
nor ( w13192 , w13191 , w11284 );
and ( w13193 , w13192 , w13367 );
and ( w13194 , w13193 , w12911 );
not ( w13195 , w13187 );
and ( w13196 , w13195 , w13194 );
nor ( w13197 , w13196 , w11099 );
and ( w13198 , w13197 , w11094 );
nor ( w13199 , w13198 , w11284 );
and ( w13200 , w13199 , w13367 );
and ( w13201 , w13200 , w12911 );
not ( w13202 , w13201 );
and ( w13203 , w13178 , w13202 );
not ( w13204 , g48 );
and ( w13205 , w13178 , w13204 );
not ( w13206 , g31 );
and ( w13207 , w13178 , w13206 );
and ( w13208 , w13207 , w13536 );
nor ( w13209 , w13205 , w13208 );
nor ( w13210 , w13209 , g47 );
not ( w13211 , g33 );
and ( w13212 , w13210 , w13211 );
and ( w13213 , w13212 , w13536 );
and ( w13214 , w13213 , w11094 );
nor ( w13215 , w13214 , w11284 );
and ( w13216 , w13215 , w13367 );
and ( w13217 , w13216 , w12911 );
not ( w13218 , w13203 );
and ( w13219 , w13218 , w13217 );
nor ( w13220 , g45 , g29 );
nor ( w13221 , w13220 , w11099 );
and ( w13222 , w13221 , w11094 );
nor ( w13223 , w13222 , w11284 );
and ( w13224 , w13223 , w13367 );
and ( w13225 , w13219 , w13224 );
nor ( w13226 , w13225 , w11186 );
nor ( w13227 , w13226 , w11284 );
and ( w13228 , w13227 , w11819 );
and ( w13229 , w13228 , w13333 );
nor ( w13230 , w13229 , w11099 );
and ( w13231 , w13230 , w11094 );
nor ( w13232 , w13231 , w11284 );
and ( w13233 , w13232 , w13367 );
and ( w13234 , w13233 , w12911 );
nor ( w13235 , g45 , w13234 );
and ( w13236 , w11703 , w11094 );
and ( w13237 , w13235 , w13236 );
and ( w13238 , w13237 , g36 );
and ( w13239 , w13238 , g11 );
nor ( w13240 , w13239 , w11284 );
and ( w13241 , w13240 , w11819 );
and ( w13242 , g45 , g29 );
and ( w13243 , w13242 , w13536 );
and ( w13244 , w13243 , w11094 );
nor ( w13245 , w13244 , w11284 );
and ( w13246 , w13245 , w13367 );
and ( w13247 , w13241 , w13246 );
and ( w13248 , w13247 , w13333 );
nor ( w13249 , w13248 , w11099 );
and ( w13250 , w13249 , w11094 );
nor ( w13251 , w13250 , w11284 );
and ( w13252 , w13251 , w13367 );
and ( w13253 , w13252 , w12911 );
nor ( w13254 , w13177 , w13253 );
and ( w13255 , w13254 , w13236 );
and ( w13256 , w13255 , w13331 );
not ( w13257 , w11186 );
and ( w13258 , w13256 , w13257 );
and ( w13259 , w13258 , w13333 );
not ( w13260 , w13259 );
and ( w13261 , w13260 , w11819 );
nor ( w13262 , w13261 , w11099 );
and ( w13263 , w13262 , w11094 );
nor ( w13264 , w13263 , w11284 );
and ( w13265 , w13264 , w13367 );
and ( w13266 , w13265 , w12911 );
not ( w13267 , w13266 );
and ( w13268 , w13161 , w13267 );
and ( w13269 , w13268 , w13492 );
not ( w13270 , w11734 );
and ( w13271 , w13269 , w13270 );
and ( w13272 , w13271 , w13563 );
nor ( w13273 , w13272 , w11284 );
and ( w13274 , w13273 , w13570 );
and ( w13275 , w13274 , w13584 );
nor ( w13276 , w13275 , w11762 );
and ( w13277 , w13157 , w13584 );
and ( w13278 , w13277 , w13367 );
and ( w13279 , w13278 , w12911 );
nor ( w13280 , g29 , w13253 );
not ( w13281 , w13280 );
and ( w13282 , w13281 , w13156 );
and ( w13283 , w13282 , w12911 );
and ( w13284 , w13279 , w13283 );
and ( w13285 , w13282 , w13084 );
and ( w13286 , w13285 , w13584 );
and ( w13287 , w13286 , w13367 );
and ( w13288 , w13287 , w12911 );
and ( w13289 , w13284 , w13288 );
nor ( w13290 , w13289 , g46 );
and ( w13291 , w13290 , w13590 );
nor ( w13292 , w13291 , w11104 );
and ( w13293 , w13292 , w13156 );
nor ( w13294 , w13293 , w11099 );
and ( w13295 , w13294 , w11094 );
nor ( w13296 , w13295 , w11284 );
and ( w13297 , w13296 , w13367 );
and ( w13298 , w13297 , w12911 );
not ( w13299 , w13276 );
and ( w13300 , w13299 , w13298 );
nor ( w13301 , w13300 , w11186 );
and ( w13302 , w13301 , w13030 );
not ( w13303 , w13302 );
and ( w13304 , w13303 , w11817 );
not ( w13305 , w13304 );
and ( w13306 , w13305 , w13236 );
not ( w13307 , w13306 );
and ( w13308 , w13307 , w13156 );
and ( w13309 , w13308 , w13084 );
not ( w13310 , w13309 );
and ( w13311 , w13310 , w11199 );
not ( w13312 , w13311 );
and ( w13313 , w13312 , w13059 );
nor ( w13314 , w13313 , w11099 );
and ( w13315 , w13314 , w11094 );
nor ( w13316 , w13315 , w11284 );
and ( w13317 , w13316 , w13367 );
and ( w13318 , w13317 , w12911 );
and ( w13319 , w13160 , w13318 );
nor ( w13320 , g43 , w11099 );
not ( w13321 , g23 );
and ( w13322 , w13320 , w13321 );
and ( w13323 , w13322 , w13492 );
and ( w13324 , w13323 , w13536 );
and ( w13325 , w13319 , w13517 );
nor ( w13326 , w13325 , w11193 );
not ( w13327 , w13326 );
and ( w13328 , w13327 , w13175 );
and ( w13329 , w13328 , w13159 );
nor ( w13330 , w13329 , w13283 );
not ( w13331 , g45 );
and ( w13332 , w13330 , w13331 );
not ( w13333 , g29 );
and ( w13334 , w13332 , w13333 );
and ( w13335 , w13334 , w13563 );
nor ( w13336 , w13335 , w11284 );
and ( w13337 , w13336 , w13570 );
and ( w13338 , w13337 , w13584 );
nor ( w13339 , w13338 , w11762 );
not ( w13340 , w13339 );
and ( w13341 , w13340 , w13298 );
nor ( w13342 , w13341 , w11186 );
and ( w13343 , w13342 , w13030 );
not ( w13344 , w13343 );
and ( w13345 , w13344 , w11817 );
not ( w13346 , w13345 );
and ( w13347 , w13346 , w13236 );
not ( w13348 , w13347 );
and ( w13349 , w13348 , w13156 );
and ( w13350 , w13349 , w13084 );
not ( w13351 , w13350 );
and ( w13352 , w13351 , w11199 );
not ( w13353 , w13352 );
and ( w13354 , w13353 , w13059 );
nor ( w13355 , w13354 , w11099 );
and ( w13356 , w13355 , w11094 );
nor ( w13357 , w13356 , w11284 );
and ( w13358 , w13357 , w13367 );
and ( w13359 , w13358 , w12911 );
and ( w13360 , w13159 , w13359 );
and ( w13361 , w13360 , w13156 );
and ( w13362 , w13361 , w13084 );
and ( w13363 , w13362 , w13367 );
and ( w13364 , w13363 , w12911 );
and ( w13365 , w13364 , w13156 );
and ( w13366 , w13365 , w12911 );
not ( w13367 , w11104 );
and ( w13368 , w13367 , w12018 );
and ( w13369 , w13584 , w13036 );
and ( w13370 , w13369 , w13084 );
and ( w13371 , w13370 , w13584 );
and ( w13372 , w13371 , w12948 );
and ( w13373 , w13372 , w12944 );
not ( w13374 , w12937 );
and ( w13375 , w13374 , w13084 );
and ( w13376 , w13375 , w13584 );
and ( w13377 , w13376 , w12948 );
and ( w13378 , w13373 , w13377 );
and ( w13379 , w13376 , w13396 );
and ( w13380 , w13379 , w13036 );
nor ( w13381 , w13380 , w11099 );
and ( w13382 , w13381 , w11094 );
not ( w13383 , w13382 );
and ( w13384 , w13383 , w13084 );
and ( w13385 , w13384 , w13584 );
and ( w13386 , w13385 , w13376 );
and ( w13387 , w13386 , w13396 );
and ( w13388 , w13387 , w13036 );
nor ( w13389 , w13388 , w11099 );
and ( w13390 , w13389 , w11094 );
not ( w13391 , w13390 );
and ( w13392 , w13391 , w13084 );
and ( w13393 , w13392 , w13584 );
and ( w13394 , w13393 , w13371 );
and ( w13395 , w13394 , w13376 );
not ( w13396 , w12935 );
and ( w13397 , w13395 , w13396 );
nor ( w13398 , w13397 , w11099 );
and ( w13399 , w13398 , w11094 );
nor ( w13400 , w13399 , w11284 );
and ( w13401 , w12948 , w13400 );
and ( w13402 , w13401 , w12944 );
and ( w13403 , w12948 , w13402 );
and ( w13404 , w13403 , w13037 );
and ( w13405 , w13084 , w12948 );
and ( w13406 , w13037 , w13405 );
and ( w13407 , w13404 , w13406 );
and ( w13408 , w13407 , w12948 );
and ( w13409 , w13408 , w13378 );
and ( w13410 , w13409 , w12944 );
and ( w13411 , w13410 , w13373 );
and ( w13412 , w13411 , w13406 );
and ( w13413 , w13412 , w12944 );
and ( w13414 , w13413 , w13377 );
and ( w13415 , w13414 , w12948 );
and ( w13416 , w13415 , w13373 );
and ( w13417 , w13416 , w13378 );
and ( w13418 , w13417 , w13373 );
and ( w13419 , w13378 , w13418 );
and ( w13420 , w13419 , w13373 );
and ( w13421 , w12948 , w13406 );
and ( w13422 , w13421 , w13037 );
and ( w13423 , w13422 , w13406 );
and ( w13424 , w13423 , w13378 );
and ( w13425 , w13424 , w12948 );
and ( w13426 , w13425 , w12944 );
and ( w13427 , w13426 , w13378 );
and ( w13428 , w13420 , w13427 );
and ( w13429 , w13428 , w13373 );
and ( w13430 , w13037 , w12944 );
and ( w13431 , w13430 , w13584 );
and ( w13432 , w13431 , w12948 );
and ( w13433 , w13432 , w13406 );
and ( w13434 , w13433 , w13570 );
and ( w13435 , w13421 , w12949 );
and ( w13436 , w13434 , w13435 );
and ( w13437 , w11186 , w13435 );
nor ( w13438 , w13437 , w12951 );
not ( w13439 , w13438 );
and ( w13440 , w13439 , w12949 );
nor ( w13441 , w13436 , w13440 );
not ( w13442 , w13441 );
and ( w13443 , w13442 , w12949 );
and ( w13444 , w13443 , w13435 );
and ( w13445 , w13444 , w13584 );
and ( w13446 , w13445 , w12948 );
and ( w13447 , w13446 , w13435 );
nor ( w13448 , w13447 , w11762 );
not ( w13449 , w13448 );
and ( w13450 , w13449 , w12948 );
and ( w13451 , w13450 , w13584 );
and ( w13452 , w13451 , w12948 );
and ( w13453 , w13452 , w13406 );
and ( w13454 , w13453 , w12948 );
and ( w13455 , w13454 , w13373 );
and ( w13456 , w13429 , w13455 );
and ( w13457 , w13456 , w13377 );
and ( w13458 , w13457 , w12948 );
and ( w13459 , w13458 , w12944 );
and ( w13460 , w13368 , w13459 );
and ( w13461 , w13366 , w13460 );
and ( w13462 , w13156 , w13460 );
and ( w13463 , w11285 , w12948 );
and ( w13464 , w13462 , w13463 );
and ( w13465 , w13461 , w13464 );
and ( w13466 , w13465 , w13460 );
and ( w13467 , w13466 , w13463 );
and ( w13468 , g45 , w13467 );
nor ( w13469 , w13468 , w12951 );
and ( w13470 , g29 , w13466 );
and ( w13471 , w13469 , w13621 );
and ( w13472 , w13041 , w13471 );
and ( w13473 , w13459 , w12948 );
not ( w13474 , g36 );
and ( w13475 , w13474 , w13473 );
nor ( w13476 , w13475 , w12951 );
not ( w13477 , g11 );
and ( w13478 , w13477 , w13459 );
and ( w13479 , w13476 , w13603 );
and ( w13480 , w13472 , w13479 );
and ( w13481 , w13480 , w13607 );
and ( w13482 , w13481 , w13556 );
and ( w13483 , w13482 , w13471 );
and ( w13484 , w13483 , w13621 );
and ( w13485 , w13584 , w13459 );
and ( w13486 , w13485 , w12948 );
not ( w13487 , w11199 );
and ( w13488 , w13487 , w13486 );
and ( w13489 , w13488 , w12949 );
nor ( w13490 , w13489 , w13440 );
and ( w13491 , w13484 , w13490 );
not ( w13492 , w9213 );
and ( w13493 , w13491 , w13492 );
not ( w13494 , w13493 );
and ( w13495 , w13494 , w12948 );
not ( w13496 , w13495 );
and ( w13497 , w13496 , w12952 );
not ( w13498 , w13497 );
and ( w13499 , w13498 , w12948 );
and ( w13500 , w13499 , w12944 );
and ( w13501 , w13500 , w13584 );
and ( w13502 , w13501 , w12948 );
not ( w13503 , w11747 );
and ( w13504 , w13502 , w13503 );
and ( w13505 , w13504 , w12949 );
and ( w13506 , w13505 , w12944 );
and ( w13507 , w13506 , w12948 );
nor ( w13508 , w13507 , w11734 );
not ( w13509 , w13508 );
and ( w13510 , w13509 , w12948 );
not ( w13511 , w9711 );
and ( w13512 , w13510 , w13511 );
not ( w13513 , w13512 );
and ( w13514 , w13513 , w12952 );
not ( w13515 , w13514 );
and ( w13516 , w13515 , w12944 );
not ( w13517 , w13324 );
and ( w13518 , w13516 , w13517 );
nor ( w13519 , w13518 , w13039 );
and ( w13520 , w13519 , w13607 );
and ( w13521 , w13520 , w13556 );
and ( w13522 , w13521 , w13479 );
and ( w13523 , w13522 , w13471 );
and ( w13524 , w13523 , w13621 );
and ( w13525 , w13524 , w13490 );
not ( w13526 , w13525 );
and ( w13527 , w13526 , w12948 );
not ( w13528 , w9108 );
and ( w13529 , w13527 , w13528 );
nor ( w13530 , w13529 , w12951 );
not ( w13531 , w13530 );
and ( w13532 , w13531 , w12948 );
not ( w13533 , w13532 );
and ( w13534 , w13533 , w12952 );
and ( w13535 , w13534 , w13607 );
not ( w13536 , w11099 );
and ( w13537 , w13535 , w13536 );
and ( w13538 , w13537 , w13607 );
and ( w13539 , w13538 , w13556 );
and ( w13540 , w13539 , w13471 );
and ( w13541 , w13540 , w13490 );
and ( w13542 , w13541 , w13471 );
and ( w13543 , w13542 , w13621 );
and ( w13544 , w13543 , w13556 );
not ( w13545 , w1853 );
and ( w13546 , w13545 , w11094 );
not ( w13547 , w13546 );
and ( w13548 , w13547 , w13084 );
and ( w13549 , w13548 , w13584 );
and ( w13550 , w13549 , w12948 );
and ( w13551 , w13544 , w13598 );
not ( w13552 , w13489 );
and ( w13553 , w13551 , w13552 );
and ( w13554 , w13553 , w13471 );
and ( w13555 , w13554 , w13490 );
not ( w13556 , w13440 );
and ( w13557 , w13555 , w13556 );
and ( w13558 , w13557 , w13471 );
and ( w13559 , w13558 , w13621 );
and ( w13560 , w13559 , w12952 );
and ( w13561 , w13560 , w13607 );
and ( w13562 , w13561 , w12952 );
not ( w13563 , w11752 );
and ( w13564 , w13562 , w13563 );
not ( w13565 , w13564 );
and ( w13566 , w13565 , w12948 );
nor ( w13567 , w13566 , w12951 );
nor ( w13568 , w13567 , w11284 );
and ( w13569 , w13568 , w12948 );
not ( w13570 , w13128 );
and ( w13571 , w13569 , w13570 );
and ( w13572 , w13571 , w13435 );
and ( w13573 , w13486 , w13435 );
and ( w13574 , w13572 , w13573 );
and ( w13575 , w13574 , w13486 );
nor ( w13576 , w13575 , w13440 );
not ( w13577 , w13576 );
and ( w13578 , w13577 , w12949 );
and ( w13579 , w13578 , w13435 );
and ( w13580 , w13459 , w13406 );
and ( w13581 , w13580 , w13037 );
and ( w13582 , w13581 , w13459 );
and ( w13583 , w13579 , w13582 );
not ( w13584 , w11284 );
and ( w13585 , w13583 , w13584 );
and ( w13586 , w13585 , w12948 );
and ( w13587 , w13586 , w13406 );
and ( w13588 , w13587 , w12948 );
nor ( w13589 , w12951 , g46 );
not ( w13590 , g9 );
and ( w13591 , w13589 , w13590 );
not ( w13592 , w13591 );
and ( w13593 , w13592 , w12944 );
and ( w13594 , w13588 , w13593 );
not ( w13595 , w13594 );
and ( w13596 , w13595 , w12952 );
and ( w13597 , w13596 , w13607 );
not ( w13598 , w13550 );
and ( w13599 , w12952 , w13598 );
and ( w13600 , w13597 , w13599 );
not ( w13601 , w13475 );
and ( w13602 , w13601 , w12952 );
not ( w13603 , w13478 );
and ( w13604 , w13602 , w13603 );
and ( w13605 , w13600 , w13604 );
and ( w13606 , w13471 , w12952 );
not ( w13607 , w12951 );
and ( w13608 , w13606 , w13607 );
and ( w13609 , w13608 , w13621 );
and ( w13610 , w13604 , w13609 );
and ( w13611 , w13610 , w13608 );
and ( w13612 , w13611 , w13604 );
and ( w13613 , w13612 , w13608 );
and ( w13614 , w13613 , w13609 );
and ( w13615 , w13614 , w13621 );
and ( w13616 , w13615 , w13604 );
and ( w13617 , w13616 , w13608 );
and ( w13618 , w13617 , w13609 );
and ( w13619 , w13618 , w13608 );
and ( w13620 , w13619 , w13609 );
not ( w13621 , w13470 );
and ( w13622 , w13620 , w13621 );
and ( w13623 , w13605 , w13622 );
and ( w13624 , w12954 , w13623 );
and ( w13625 , w13627 , w12944 );
and ( w13626 , w13625 , w13463 );
not ( w13627 , w13624 );
and ( w13628 , w13626 , w13627 );
and ( w13629 , w13628 , w13461 );
and ( w13630 , w13629 , w13465 );
and ( t_3 , w13630 , w13461 );

endmodule
