module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 ; 
output g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
n2870 , n2871 , n2872 , n2873 ; 
wire t_0 , t_1 , t_2 , t_3 , t_4 , t_5 , t_6 , t_7 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( g136 , n137 ); 
buf ( g137 , n138 ); 
buf ( g138 , n139 ); 
buf ( g139 , n140 ); 
buf ( g140 , n141 ); 
buf ( g141 , n142 ); 
buf ( g142 , n143 ); 
buf ( g143 , n144 ); 
buf ( g144 , n145 ); 
buf ( g145 , n146 ); 
buf ( g146 , n147 ); 
buf ( g147 , n148 ); 
buf ( g148 , n149 ); 
buf ( g149 , n150 ); 
buf ( g150 , n151 ); 
buf ( g151 , n152 ); 
buf ( g152 , n153 ); 
buf ( g153 , n154 ); 
buf ( g154 , n155 ); 
buf ( g155 , n156 ); 
buf ( g156 , n157 ); 
buf ( g157 , n158 ); 
buf ( g158 , n159 ); 
buf ( g159 , n160 ); 
buf ( g160 , n161 ); 
buf ( g161 , n162 ); 
buf ( g162 , n163 ); 
buf ( g163 , n164 ); 
buf ( g164 , n165 ); 
buf ( g165 , n166 ); 
buf ( g166 , n167 ); 
buf ( n137 , n2320 ); 
buf ( n138 , n1301 ); 
buf ( n139 , n1377 ); 
buf ( n140 , n633 ); 
buf ( n141 , n713 ); 
buf ( n142 , n2873 ); 
buf ( n143 , n1608 ); 
buf ( n144 , n1690 ); 
buf ( n145 , n718 ); 
buf ( n146 , n1696 ); 
buf ( n147 , n2722 ); 
buf ( n148 , n2517 ); 
buf ( n149 , n2180 ); 
buf ( n150 , n1751 ); 
buf ( n151 , n2229 ); 
buf ( n152 , n2866 ); 
buf ( n153 , n1823 ); 
buf ( n154 , n775 ); 
buf ( n155 , n1005 ); 
buf ( n156 , n2614 ); 
buf ( n157 , n2782 ); 
buf ( n158 , n1880 ); 
buf ( n159 , n2108 ); 
buf ( n160 , n1083 ); 
buf ( n161 , n2816 ); 
buf ( n162 , n2609 ); 
buf ( n163 , n2547 ); 
buf ( n164 , n2668 ); 
buf ( n165 , n404 ); 
buf ( n166 , n2185 ); 
buf ( n167 , n1818 ); 
not ( n170 , n132 ); 
not ( n171 , n170 ); 
and ( n172 , n64 , n63 ); 
not ( n173 , n64 ); 
not ( n174 , n63 ); 
and ( n175 , n173 , n174 ); 
nor ( n176 , n172 , n175 ); 
not ( n177 , n176 ); 
buf ( n178 , n177 ); 
not ( n179 , n178 ); 
not ( n180 , n179 ); 
xor ( n181 , n71 , n72 ); 
buf ( n182 , n181 ); 
not ( n183 , n182 ); 
and ( n184 , n70 , n69 ); 
not ( n185 , n70 ); 
not ( n186 , n69 ); 
and ( n187 , n185 , n186 ); 
nor ( n188 , n184 , n187 ); 
not ( n189 , n188 ); 
not ( n190 , n189 ); 
and ( n191 , n66 , n65 ); 
not ( n192 , n66 ); 
not ( n193 , n65 ); 
and ( n194 , n192 , n193 ); 
nor ( n195 , n191 , n194 ); 
not ( n196 , n67 ); 
and ( n197 , n68 , n196 ); 
not ( n198 , n68 ); 
and ( n199 , n198 , n67 ); 
nor ( n200 , n197 , n199 ); 
not ( n201 , n200 ); 
nand ( n202 , n190 , n195 , n201 ); 
not ( n203 , n202 ); 
nand ( n204 , n183 , n203 ); 
and ( n205 , n62 , n61 ); 
not ( n206 , n62 ); 
not ( n207 , n61 ); 
and ( n208 , n206 , n207 ); 
nor ( n209 , n205 , n208 ); 
buf ( n210 , n209 ); 
not ( n211 , n210 ); 
nor ( n212 , n204 , n211 ); 
nand ( n213 , n180 , n212 ); 
buf ( n214 , n188 ); 
nand ( n215 , n214 , n195 ); 
not ( n216 , n200 ); 
nor ( n217 , n215 , n216 ); 
nand ( n218 , n182 , n217 ); 
not ( n219 , n218 ); 
not ( n220 , n209 ); 
not ( n221 , n220 ); 
buf ( n222 , n221 ); 
nand ( n223 , n219 , n222 , n180 ); 
and ( n224 , n213 , n223 ); 
not ( n225 , n178 ); 
not ( n226 , n189 ); 
xor ( n227 , n66 , n65 ); 
not ( n228 , n227 ); 
nand ( n229 , n226 , n216 , n228 ); 
not ( n230 , n182 ); 
nor ( n231 , n229 , n230 ); 
nand ( n232 , n225 , n222 , n231 ); 
nor ( n233 , n182 , n229 ); 
nand ( n234 , n180 , n222 , n233 ); 
and ( n235 , n232 , n234 ); 
not ( n236 , n225 ); 
not ( n237 , n209 ); 
not ( n238 , n237 ); 
not ( n239 , n195 ); 
buf ( n240 , n200 ); 
nand ( n241 , n239 , n226 , n240 ); 
nor ( n242 , n182 , n241 ); 
nand ( n243 , n238 , n242 ); 
nor ( n244 , n236 , n243 ); 
not ( n245 , n244 ); 
not ( n246 , n178 ); 
buf ( n247 , n220 ); 
not ( n248 , n247 ); 
buf ( n249 , n181 ); 
not ( n250 , n249 ); 
not ( n251 , n250 ); 
not ( n252 , n214 ); 
nand ( n253 , n252 , n216 , n227 ); 
not ( n254 , n253 ); 
nand ( n255 , n251 , n254 ); 
not ( n256 , n255 ); 
nand ( n257 , n246 , n248 , n256 ); 
not ( n258 , n257 ); 
buf ( n259 , n177 ); 
buf ( n260 , n259 ); 
not ( n261 , n260 ); 
nor ( n262 , n250 , n202 ); 
nand ( n263 , n221 , n262 ); 
not ( n264 , n263 ); 
not ( n265 , n264 ); 
or ( n266 , n261 , n265 ); 
not ( n267 , n217 ); 
nor ( n268 , n251 , n267 ); 
not ( n269 , n178 ); 
nand ( n270 , n268 , n238 , n269 ); 
nand ( n271 , n266 , n270 ); 
nor ( n272 , n258 , n271 ); 
nand ( n273 , n224 , n235 , n245 , n272 ); 
not ( n274 , n259 ); 
nor ( n275 , n253 , n182 ); 
nand ( n276 , n274 , n211 , n275 ); 
not ( n277 , n178 ); 
not ( n278 , n195 ); 
and ( n279 , n200 , n278 , n189 ); 
and ( n280 , n220 , n182 , n279 ); 
nand ( n281 , n277 , n280 ); 
and ( n282 , n276 , n281 ); 
not ( n283 , n260 ); 
not ( n284 , n210 ); 
and ( n285 , n284 , n242 ); 
and ( n286 , n283 , n285 ); 
not ( n287 , n231 ); 
nor ( n288 , n209 , n176 ); 
not ( n289 , n288 ); 
not ( n290 , n289 ); 
not ( n291 , n290 ); 
nor ( n292 , n287 , n291 ); 
nor ( n293 , n286 , n292 ); 
and ( n294 , n260 , n285 ); 
not ( n295 , n260 ); 
not ( n296 , n240 ); 
nor ( n297 , n227 , n214 ); 
nand ( n298 , n296 , n297 ); 
not ( n299 , n182 ); 
nor ( n300 , n298 , n299 ); 
and ( n301 , n247 , n300 ); 
and ( n302 , n295 , n301 ); 
nor ( n303 , n294 , n302 ); 
nand ( n304 , n282 , n293 , n303 ); 
not ( n305 , n304 ); 
not ( n306 , n220 ); 
buf ( n307 , n189 ); 
not ( n308 , n228 ); 
nand ( n309 , n307 , n308 , n240 ); 
nor ( n310 , n309 , n299 ); 
nand ( n311 , n306 , n310 ); 
nor ( n312 , n311 , n225 ); 
nand ( n313 , n178 , n238 , n300 ); 
not ( n314 , n313 ); 
nor ( n315 , n312 , n314 ); 
nand ( n316 , n275 , n306 ); 
not ( n317 , n269 ); 
nor ( n318 , n316 , n317 ); 
not ( n319 , n279 ); 
not ( n320 , n249 ); 
nor ( n321 , n319 , n320 ); 
nand ( n322 , n238 , n321 ); 
nor ( n323 , n260 , n322 ); 
nor ( n324 , n318 , n323 ); 
nand ( n325 , n179 , n211 , n262 ); 
nor ( n326 , n177 , n249 ); 
not ( n327 , n237 ); 
nand ( n328 , n326 , n327 , n279 ); 
nand ( n329 , n325 , n328 ); 
nand ( n330 , n274 , n211 , n233 ); 
nor ( n331 , n182 , n298 ); 
nand ( n332 , n274 , n238 , n331 ); 
nand ( n333 , n330 , n332 ); 
nor ( n334 , n329 , n333 ); 
and ( n335 , n315 , n324 , n334 ); 
not ( n336 , n296 ); 
not ( n337 , n336 ); 
not ( n338 , n337 ); 
not ( n339 , n338 ); 
not ( n340 , n221 ); 
not ( n341 , n308 ); 
nand ( n342 , n214 , n181 ); 
or ( n343 , n341 , n177 , n342 ); 
not ( n344 , n189 ); 
nor ( n345 , n344 , n181 ); 
not ( n346 , n227 ); 
nand ( n347 , n345 , n177 , n346 ); 
nand ( n348 , n343 , n347 ); 
not ( n349 , n348 ); 
or ( n350 , n340 , n349 ); 
not ( n351 , n342 ); 
nand ( n352 , n351 , n341 , n288 ); 
nand ( n353 , n350 , n352 ); 
not ( n354 , n353 ); 
or ( n355 , n339 , n354 ); 
not ( n356 , n341 ); 
not ( n357 , n356 ); 
not ( n358 , n289 ); 
nand ( n359 , n357 , n337 , n358 , n345 ); 
nand ( n360 , n355 , n359 ); 
not ( n361 , n360 ); 
nor ( n362 , n222 , n255 ); 
nand ( n363 , n260 , n362 ); 
not ( n364 , n260 ); 
nor ( n365 , n309 , n182 ); 
nand ( n366 , n365 , n247 ); 
not ( n367 , n366 ); 
nand ( n368 , n364 , n367 ); 
nand ( n369 , n361 , n363 , n368 ); 
nor ( n370 , n366 , n246 ); 
not ( n371 , n370 ); 
nand ( n372 , n280 , n260 ); 
nand ( n373 , n371 , n372 ); 
nor ( n374 , n369 , n373 ); 
nor ( n375 , n204 , n327 ); 
not ( n376 , n375 ); 
nor ( n377 , n283 , n376 ); 
not ( n378 , n377 ); 
nor ( n379 , n218 , n306 ); 
nand ( n380 , n260 , n379 ); 
and ( n381 , n378 , n380 ); 
nand ( n382 , n305 , n335 , n374 , n381 ); 
nor ( n383 , n273 , n382 ); 
not ( n384 , n383 ); 
or ( n385 , n171 , n384 ); 
not ( n386 , n17 ); 
not ( n387 , n18 ); 
not ( n388 , n3 ); 
not ( n389 , n19 ); 
or ( n390 , n386 , n387 , n388 , n389 ); 
buf ( n391 , n390 ); 
nand ( n392 , n385 , n391 ); 
not ( n393 , n273 ); 
not ( n394 , n374 ); 
not ( n395 , n304 ); 
nand ( n396 , n395 , n381 ); 
nor ( n397 , n394 , n396 ); 
and ( n398 , n393 , n335 , n397 ); 
nor ( n399 , n398 , n170 ); 
or ( n400 , n392 , n399 ); 
not ( n401 , n133 ); 
buf ( n402 , n390 ); 
or ( n403 , n401 , n402 ); 
nand ( n404 , n400 , n403 ); 
not ( n405 , n39 ); 
not ( n406 , n405 ); 
xor ( n407 , n40 , n41 ); 
not ( n408 , n407 ); 
buf ( n409 , n408 ); 
and ( n410 , n46 , n47 ); 
not ( n411 , n46 ); 
not ( n412 , n47 ); 
and ( n413 , n411 , n412 ); 
nor ( n414 , n410 , n413 ); 
buf ( n415 , n414 ); 
and ( n416 , n42 , n43 ); 
not ( n417 , n42 ); 
not ( n418 , n43 ); 
and ( n419 , n417 , n418 ); 
nor ( n420 , n416 , n419 ); 
not ( n421 , n420 ); 
not ( n422 , n421 ); 
xor ( n423 , n50 , n51 ); 
and ( n424 , n415 , n422 , n423 ); 
and ( n425 , n48 , n49 ); 
not ( n426 , n48 ); 
not ( n427 , n49 ); 
and ( n428 , n426 , n427 ); 
nor ( n429 , n425 , n428 ); 
not ( n430 , n429 ); 
nand ( n431 , n424 , n430 ); 
not ( n432 , n44 ); 
not ( n433 , n45 ); 
not ( n434 , n433 ); 
or ( n435 , n432 , n434 ); 
not ( n436 , n44 ); 
nand ( n437 , n45 , n436 ); 
nand ( n438 , n435 , n437 ); 
not ( n439 , n438 ); 
not ( n440 , n439 ); 
nor ( n441 , n431 , n440 ); 
nand ( n442 , n409 , n441 ); 
buf ( n443 , n438 ); 
not ( n444 , n443 ); 
not ( n445 , n429 ); 
not ( n446 , n445 ); 
buf ( n447 , n408 ); 
not ( n448 , n414 ); 
and ( n449 , n448 , n422 , n423 ); 
nand ( n450 , n444 , n446 , n447 , n449 ); 
nand ( n451 , n442 , n450 ); 
buf ( n452 , n407 ); 
buf ( n453 , n439 ); 
and ( n454 , n48 , n427 ); 
not ( n455 , n48 ); 
and ( n456 , n455 , n49 ); 
or ( n457 , n454 , n456 ); 
not ( n458 , n457 ); 
and ( n459 , n50 , n51 ); 
not ( n460 , n50 ); 
not ( n461 , n51 ); 
and ( n462 , n460 , n461 ); 
nor ( n463 , n459 , n462 ); 
not ( n464 , n463 ); 
not ( n465 , n420 ); 
and ( n466 , n464 , n465 , n414 ); 
nand ( n467 , n458 , n466 ); 
not ( n468 , n467 ); 
nand ( n469 , n452 , n453 , n468 ); 
not ( n470 , n469 ); 
not ( n471 , n470 ); 
not ( n472 , n414 ); 
not ( n473 , n421 ); 
nor ( n474 , n473 , n463 ); 
and ( n475 , n472 , n474 ); 
not ( n476 , n475 ); 
nor ( n477 , n446 , n476 ); 
not ( n478 , n447 ); 
nand ( n479 , n477 , n444 , n478 ); 
nand ( n480 , n471 , n479 ); 
not ( n481 , n480 ); 
not ( n482 , n407 ); 
buf ( n483 , n482 ); 
not ( n484 , n472 ); 
not ( n485 , n420 ); 
nand ( n486 , n485 , n463 ); 
not ( n487 , n486 ); 
nand ( n488 , n430 , n484 , n487 ); 
nor ( n489 , n488 , n440 ); 
nand ( n490 , n483 , n489 ); 
not ( n491 , n438 ); 
not ( n492 , n415 ); 
and ( n493 , n491 , n430 , n492 , n487 ); 
nand ( n494 , n483 , n493 ); 
nand ( n495 , n481 , n490 , n494 ); 
nor ( n496 , n451 , n495 ); 
not ( n497 , n447 ); 
not ( n498 , n463 ); 
not ( n499 , n465 ); 
not ( n500 , n414 ); 
nand ( n501 , n498 , n499 , n500 ); 
not ( n502 , n501 ); 
not ( n503 , n445 ); 
nand ( n504 , n502 , n503 ); 
nor ( n505 , n453 , n504 ); 
nand ( n506 , n497 , n505 ); 
not ( n507 , n506 ); 
not ( n508 , n409 ); 
not ( n509 , n508 ); 
buf ( n510 , n445 ); 
nand ( n511 , n510 , n449 ); 
nor ( n512 , n453 , n511 ); 
not ( n513 , n512 ); 
or ( n514 , n509 , n513 ); 
not ( n515 , n447 ); 
not ( n516 , n491 ); 
not ( n517 , n431 ); 
nand ( n518 , n515 , n516 , n517 ); 
nand ( n519 , n514 , n518 ); 
nor ( n520 , n507 , n519 ); 
buf ( n521 , n408 ); 
not ( n522 , n521 ); 
not ( n523 , n445 ); 
and ( n524 , n443 , n523 , n466 ); 
nand ( n525 , n522 , n524 ); 
not ( n526 , n522 ); 
nand ( n527 , n430 , n492 , n487 ); 
nor ( n528 , n453 , n527 ); 
not ( n529 , n528 ); 
nor ( n530 , n526 , n529 ); 
buf ( n531 , n499 ); 
nand ( n532 , n531 , n415 , n457 , n423 ); 
nor ( n533 , n453 , n532 ); 
nand ( n534 , n483 , n533 ); 
not ( n535 , n452 ); 
nand ( n536 , n535 , n512 ); 
nand ( n537 , n496 , n520 , t_2 ); 
nor ( n538 , n407 , n438 ); 
not ( n539 , n423 ); 
nand ( n540 , n539 , n531 , n415 ); 
nor ( n541 , n540 , n510 ); 
nand ( n542 , n538 , n541 ); 
and ( n543 , n475 , n523 , n491 ); 
nand ( n544 , n543 , n409 ); 
and ( n545 , n542 , n544 ); 
not ( n546 , n415 ); 
nor ( n547 , n546 , n486 ); 
nand ( n548 , n523 , n443 , n547 ); 
nor ( n549 , n483 , n548 ); 
not ( n550 , n549 ); 
nand ( n551 , n545 , n550 ); 
not ( n552 , n472 ); 
not ( n553 , n552 ); 
not ( n554 , n523 ); 
nor ( n555 , n553 , n554 ); 
not ( n556 , n422 ); 
not ( n557 , n556 ); 
buf ( n558 , n440 ); 
not ( n559 , n558 ); 
not ( n560 , n423 ); 
nand ( n561 , n560 , n407 ); 
not ( n562 , n561 ); 
nand ( n563 , n555 , n557 , n559 , n562 ); 
not ( n564 , n502 ); 
not ( n565 , n564 ); 
not ( n566 , n523 ); 
nand ( n567 , n565 , n566 , n453 ); 
not ( n568 , n567 ); 
nand ( n569 , n526 , n568 ); 
nand ( n570 , n457 , n423 ); 
nor ( n571 , n492 , n438 , n570 ); 
not ( n572 , n571 ); 
nor ( n573 , n457 , n423 ); 
not ( n574 , n573 ); 
nand ( n575 , n574 , n570 ); 
nand ( n576 , n553 , n440 , n575 ); 
nand ( n577 , n572 , n576 ); 
buf ( n578 , n521 ); 
nand ( n579 , n577 , n578 , n556 ); 
nand ( n580 , n563 , n569 , n579 ); 
nor ( n581 , n551 , n580 ); 
not ( n582 , n578 ); 
not ( n583 , n523 ); 
not ( n584 , n540 ); 
nand ( n585 , n583 , n584 ); 
nor ( n586 , n585 , n516 ); 
nand ( n587 , n582 , n586 ); 
nand ( n588 , n582 , n543 ); 
and ( n589 , n587 , n588 ); 
not ( n590 , n585 ); 
nand ( n591 , n535 , n558 , n590 ); 
not ( n592 , n511 ); 
nand ( n593 , n497 , n559 , n592 ); 
and ( n594 , n591 , n593 ); 
nand ( n595 , n478 , n489 ); 
not ( n596 , n595 ); 
nand ( n597 , n409 , n505 ); 
not ( n598 , n597 ); 
nor ( n599 , n596 , n598 ); 
nand ( n600 , n409 , n524 ); 
not ( n601 , n600 ); 
not ( n602 , n564 ); 
not ( n603 , n521 ); 
nand ( n604 , n602 , n603 , n440 , n554 ); 
not ( n605 , n604 ); 
nor ( n606 , n601 , n605 ); 
nor ( n607 , n453 , n467 ); 
nand ( n608 , n409 , n607 ); 
not ( n609 , n608 ); 
nand ( n610 , n452 , n446 , n491 , n449 ); 
not ( n611 , n610 ); 
nor ( n612 , n609 , n611 ); 
nand ( n613 , n599 , n606 , n612 ); 
not ( n614 , n613 ); 
nand ( n615 , n581 , n589 , n594 , n614 ); 
nor ( n616 , n537 , n615 ); 
not ( n617 , n616 ); 
or ( n618 , n406 , n617 ); 
not ( n619 , n391 ); 
nand ( n620 , n618 , n619 ); 
not ( n621 , n537 ); 
not ( n622 , n581 ); 
nand ( n623 , n594 , n599 , n606 , n612 ); 
nor ( n624 , n622 , n623 ); 
and ( n625 , n621 , n589 , n624 ); 
nor ( n626 , n625 , n405 ); 
or ( n627 , n620 , n626 ); 
and ( n628 , n38 , n388 ); 
and ( n629 , n1 , n3 ); 
nor ( n630 , n628 , n629 ); 
not ( n631 , n391 ); 
or ( n632 , n630 , n631 ); 
nand ( n633 , n627 , n632 ); 
and ( n634 , n52 , n388 ); 
and ( n635 , n3 , n20 ); 
nor ( n636 , n634 , n635 ); 
and ( n637 , n391 , n636 ); 
not ( n638 , n391 ); 
nand ( n639 , n526 , n586 ); 
nand ( n640 , n639 , n569 ); 
not ( n641 , n553 ); 
and ( n642 , n45 , n44 ); 
not ( n643 , n45 ); 
and ( n644 , n643 , n436 ); 
nor ( n645 , n642 , n644 ); 
not ( n646 , n645 ); 
nand ( n647 , n556 , n646 ); 
not ( n648 , n423 ); 
nor ( n649 , n648 , n407 ); 
not ( n650 , n649 ); 
nand ( n651 , n650 , n561 ); 
or ( n652 , n554 , n647 , n651 ); 
nand ( n653 , n531 , n645 ); 
not ( n654 , n653 ); 
nand ( n655 , n566 , n654 , n651 ); 
nand ( n656 , n652 , n655 ); 
nand ( n657 , n641 , n656 ); 
nand ( n658 , n497 , n533 ); 
nor ( n659 , n552 , n486 ); 
and ( n660 , n407 , n457 ); 
nand ( n661 , n659 , n440 , n660 ); 
nand ( n662 , n657 , n658 , n661 ); 
nor ( n663 , n640 , n662 ); 
not ( n664 , n450 ); 
not ( n665 , n664 ); 
not ( n666 , n578 ); 
nand ( n667 , n666 , n568 ); 
nand ( n668 , n665 , n667 ); 
not ( n669 , n482 ); 
not ( n670 , n504 ); 
nand ( n671 , n669 , n670 , n453 ); 
not ( n672 , n671 ); 
nor ( n673 , n672 , n470 ); 
nand ( n674 , n673 , n490 , n494 ); 
nor ( n675 , n668 , n674 ); 
and ( n676 , n663 , n545 , n675 ); 
not ( n677 , n604 ); 
not ( n678 , n521 ); 
nor ( n679 , n678 , n548 ); 
nor ( n680 , n677 , n679 ); 
not ( n681 , n518 ); 
nor ( n682 , n681 , n530 ); 
not ( n683 , n525 ); 
not ( n684 , n536 ); 
nor ( n685 , n683 , n684 ); 
and ( n686 , t_0 , n680 , n682 , n685 ); 
not ( n687 , n532 ); 
nand ( n688 , n687 , n444 ); 
not ( n689 , n688 ); 
nand ( n690 , n689 , n578 ); 
not ( n691 , n690 ); 
nand ( n692 , n508 , n493 ); 
not ( n693 , n692 ); 
nor ( n694 , n691 , n693 ); 
not ( n695 , n441 ); 
nor ( n696 , n695 , n578 ); 
nor ( n697 , n696 , n611 ); 
not ( n698 , n591 ); 
nand ( n699 , n535 , n516 , n541 ); 
not ( n700 , n699 ); 
nor ( n701 , n698 , n700 ); 
nor ( n702 , n566 , n476 ); 
and ( n703 , n483 , n558 , n702 ); 
not ( n704 , n608 ); 
nor ( n705 , n703 , n704 ); 
and ( n706 , n694 , n697 , n701 , n705 ); 
nand ( n707 , n676 , n686 , n706 ); 
not ( n708 , n53 ); 
and ( n709 , n707 , n708 ); 
and ( n710 , t_5 , n53 ); 
nor ( n711 , n709 , n710 ); 
and ( n712 , n638 , n711 ); 
nor ( n713 , n637 , n712 ); 
not ( n714 , n73 ); 
and ( n715 , n631 , n714 ); 
not ( n716 , n631 ); 
and ( n717 , n716 , n711 ); 
nor ( n718 , n715 , n717 ); 
not ( n719 , n111 ); 
not ( n720 , n719 ); 
not ( n721 , n466 ); 
nor ( n722 , n510 , n721 ); 
nand ( n723 , n722 , n453 , n452 ); 
and ( n724 , n671 , n723 ); 
nand ( n725 , n724 , n490 , n479 ); 
nor ( n726 , t_7 , n725 ); 
not ( n727 , n478 ); 
not ( n728 , n607 ); 
or ( n729 , n727 , n728 ); 
nand ( n730 , n729 , n604 ); 
nor ( n731 , n681 , n730 ); 
not ( n732 , n661 ); 
nor ( n733 , n732 , n679 ); 
nand ( n734 , n409 , n528 ); 
and ( n735 , n534 , n733 , n536 , n734 ); 
and ( n736 , n726 , n731 , n735 ); 
not ( n737 , n736 ); 
and ( n738 , n699 , n610 ); 
not ( n739 , n608 ); 
nor ( n740 , n688 , n483 ); 
nor ( n741 , n739 , n740 ); 
and ( n742 , n597 , n600 ); 
nand ( n743 , n738 , n741 , n742 ); 
not ( n744 , n743 ); 
not ( n745 , n549 ); 
not ( n746 , n423 ); 
nand ( n747 , n746 , n552 , n654 ); 
nor ( n748 , n746 , n484 ); 
nand ( n749 , n653 , n647 ); 
nand ( n750 , n748 , n749 ); 
nand ( n751 , n747 , n750 ); 
not ( n752 , n554 ); 
nand ( n753 , n751 , n497 , n752 ); 
nand ( n754 , n745 , n569 , n753 ); 
not ( n755 , n647 ); 
nand ( n756 , n755 , n641 , n409 , n573 ); 
nand ( n757 , n756 , n639 , n544 ); 
nor ( n758 , n754 , n757 ); 
buf ( n759 , n694 ); 
nand ( n760 , n744 , n758 , n759 , t_4 ); 
nor ( n761 , n737 , n760 ); 
not ( n762 , n761 ); 
or ( n763 , n720 , n762 ); 
nand ( n764 , n763 , n402 ); 
buf ( n765 , n736 ); 
not ( n766 , n758 ); 
nand ( n767 , t_3 , n738 , n741 , n742 ); 
nor ( n768 , n766 , n767 ); 
buf ( n769 , n759 ); 
and ( n770 , n765 , n768 , n769 ); 
nor ( n771 , n770 , n719 ); 
or ( n772 , n764 , n771 ); 
not ( n773 , n112 ); 
or ( n774 , n773 , n402 ); 
nand ( n775 , n772 , n774 ); 
xor ( n776 , n6 , n105 ); 
not ( n777 , n776 ); 
not ( n778 , n777 ); 
not ( n779 , n778 ); 
not ( n780 , n779 ); 
and ( n781 , n98 , n99 ); 
not ( n782 , n98 ); 
not ( n783 , n99 ); 
and ( n784 , n782 , n783 ); 
nor ( n785 , n781 , n784 ); 
buf ( n786 , n785 ); 
not ( n787 , n786 ); 
not ( n788 , n787 ); 
xor ( n789 , n101 , n102 ); 
buf ( n790 , n789 ); 
not ( n791 , n790 ); 
and ( n792 , n62 , n103 ); 
not ( n793 , n62 ); 
not ( n794 , n103 ); 
and ( n795 , n793 , n794 ); 
nor ( n796 , n792 , n795 ); 
buf ( n797 , n796 ); 
not ( n798 , n104 ); 
not ( n799 , n64 ); 
not ( n800 , n799 ); 
or ( n801 , n798 , n800 ); 
not ( n802 , n104 ); 
nand ( n803 , n64 , n802 ); 
nand ( n804 , n801 , n803 ); 
nand ( n805 , n797 , n804 ); 
not ( n806 , n805 ); 
nand ( n807 , n788 , n791 , n806 ); 
xor ( n808 , n8 , n100 ); 
not ( n809 , n808 ); 
buf ( n810 , n809 ); 
not ( n811 , n810 ); 
nor ( n812 , n807 , n811 ); 
nand ( n813 , n780 , n812 ); 
nor ( n814 , n808 , n776 ); 
not ( n815 , n786 ); 
not ( n816 , n796 ); 
nor ( n817 , n816 , n804 ); 
nand ( n818 , n815 , n817 ); 
not ( n819 , n789 ); 
not ( n820 , n819 ); 
nor ( n821 , n818 , n820 ); 
nand ( n822 , n814 , n821 ); 
nor ( n823 , n804 , n796 ); 
not ( n824 , n785 ); 
and ( n825 , n823 , n824 ); 
not ( n826 , n789 ); 
nand ( n827 , n825 , n826 ); 
not ( n828 , n827 ); 
nor ( n829 , n808 , n776 ); 
nand ( n830 , n828 , n829 ); 
and ( n831 , n822 , n830 ); 
and ( n832 , n813 , n831 ); 
not ( n833 , n778 ); 
not ( n834 , n833 ); 
not ( n835 , n834 ); 
buf ( n836 , n808 ); 
not ( n837 , n836 ); 
buf ( n838 , n789 ); 
not ( n839 , n838 ); 
nor ( n840 , n818 , n839 ); 
nand ( n841 , n837 , n840 ); 
not ( n842 , n841 ); 
not ( n843 , n842 ); 
or ( n844 , n835 , n843 ); 
not ( n845 , n777 ); 
buf ( n846 , n845 ); 
not ( n847 , n804 ); 
not ( n848 , n824 ); 
not ( n849 , n797 ); 
not ( n850 , n849 ); 
nand ( n851 , n847 , n848 , n850 , n838 ); 
not ( n852 , n810 ); 
nor ( n853 , n851 , n852 ); 
nand ( n854 , n846 , n853 ); 
nand ( n855 , n844 , n854 ); 
not ( n856 , n855 ); 
buf ( n857 , n778 ); 
not ( n858 , n852 ); 
not ( n859 , n848 ); 
nand ( n860 , n839 , n859 , n806 ); 
not ( n861 , n860 ); 
nand ( n862 , n857 , n858 , n861 ); 
nand ( n863 , n810 , n777 ); 
not ( n864 , n796 ); 
nand ( n865 , n864 , n804 ); 
not ( n866 , n865 ); 
and ( n867 , n826 , n787 , n866 ); 
not ( n868 , n867 ); 
nor ( n869 , n863 , n868 ); 
not ( n870 , n869 ); 
and ( n871 , n862 , n870 ); 
buf ( n872 , n776 ); 
not ( n873 , n872 ); 
nand ( n874 , n873 , n836 , n821 ); 
not ( n875 , n874 ); 
not ( n876 , n875 ); 
nand ( n877 , n866 , n848 ); 
not ( n878 , n877 ); 
not ( n879 , n820 ); 
nand ( n880 , n878 , n879 ); 
not ( n881 , n880 ); 
not ( n882 , n776 ); 
buf ( n883 , n882 ); 
not ( n884 , n883 ); 
not ( n885 , n836 ); 
not ( n886 , n885 ); 
nand ( n887 , n881 , n884 , n886 ); 
nand ( n888 , n876 , n887 ); 
not ( n889 , n873 ); 
not ( n890 , n790 ); 
not ( n891 , n817 ); 
nor ( n892 , n891 , n787 ); 
nand ( n893 , n890 , n892 ); 
not ( n894 , n893 ); 
nand ( n895 , n889 , n811 , n894 ); 
not ( n896 , n847 ); 
not ( n897 , n786 ); 
or ( n898 , n896 , n897 , n819 ); 
nand ( n899 , n896 , n897 , n826 ); 
nand ( n900 , n898 , n899 ); 
not ( n901 , n777 ); 
not ( n902 , n808 ); 
nor ( n903 , n849 , n902 ); 
not ( n904 , n903 ); 
not ( n905 , n808 ); 
nand ( n906 , n905 , n849 ); 
nand ( n907 , n904 , n906 ); 
nand ( n908 , n900 , n901 , n907 ); 
nand ( n909 , n895 , n908 ); 
nor ( n910 , n888 , n909 ); 
nand ( n911 , n832 , n856 , n871 , n910 ); 
not ( n912 , n889 ); 
not ( n913 , n912 ); 
not ( n914 , n836 ); 
nor ( n915 , n807 , n914 ); 
not ( n916 , n915 ); 
or ( n917 , n913 , n916 ); 
not ( n918 , n836 ); 
not ( n919 , n918 ); 
nand ( n920 , n919 , n833 , n861 ); 
nand ( n921 , n917 , n920 ); 
not ( n922 , n921 ); 
buf ( n923 , n836 ); 
nor ( n924 , n804 , n797 ); 
and ( n925 , n786 , n924 ); 
not ( n926 , n925 ); 
nor ( n927 , n879 , n926 ); 
nand ( n928 , n779 , n923 , n927 ); 
nand ( n929 , n839 , n925 ); 
not ( n930 , n929 ); 
not ( n931 , n845 ); 
nand ( n932 , n930 , n858 , n931 ); 
and ( n933 , n928 , n932 ); 
nor ( n934 , n787 , n805 ); 
nand ( n935 , n790 , n934 ); 
not ( n936 , n935 ); 
nand ( n937 , n884 , n886 , n936 ); 
not ( n938 , n937 ); 
not ( n939 , n885 ); 
not ( n940 , n877 ); 
nand ( n941 , n940 , n790 ); 
not ( n942 , n941 ); 
nand ( n943 , n939 , n942 , n779 ); 
not ( n944 , n943 ); 
nor ( n945 , n938 , n944 ); 
not ( n946 , n805 ); 
nand ( n947 , n946 , n790 , n859 ); 
not ( n948 , n947 ); 
nand ( n949 , n857 , n886 , n948 ); 
not ( n950 , n941 ); 
not ( n951 , n852 ); 
nand ( n952 , n950 , n857 , n951 ); 
and ( n953 , n949 , n952 ); 
nand ( n954 , n922 , n933 , n945 , n953 ); 
nor ( n955 , n911 , n954 ); 
not ( n956 , n825 ); 
not ( n957 , n790 ); 
nor ( n958 , n956 , n957 ); 
not ( n959 , n958 ); 
nor ( n960 , n959 , n914 ); 
not ( n961 , n960 ); 
not ( n962 , n901 ); 
not ( n963 , n962 ); 
nor ( n964 , n961 , n963 ); 
not ( n965 , n819 ); 
nand ( n966 , n859 , n965 , n866 ); 
nor ( n967 , n951 , n966 ); 
not ( n968 , n967 ); 
not ( n969 , n883 ); 
not ( n970 , n969 ); 
nor ( n971 , n968 , n970 ); 
nor ( n972 , n964 , n971 ); 
nand ( n973 , n780 , n960 ); 
nor ( n974 , n811 , n893 ); 
nand ( n975 , n780 , n974 ); 
and ( n976 , n973 , n975 ); 
not ( n977 , n812 ); 
nor ( n978 , n977 , n963 ); 
nor ( n979 , n846 , n841 ); 
nor ( n980 , n978 , n979 ); 
and ( n981 , n972 , n976 , n980 ); 
not ( n982 , n851 ); 
nand ( n983 , n982 , n811 , n883 ); 
not ( n984 , n983 ); 
nor ( n985 , n827 , n885 ); 
nand ( n986 , n985 , n884 ); 
not ( n987 , n986 ); 
nor ( n988 , n984 , n987 ); 
not ( n989 , n966 ); 
and ( n990 , n833 , n858 , n989 ); 
nor ( n991 , n811 , n947 ); 
nand ( n992 , n962 , n991 ); 
not ( n993 , n992 ); 
nor ( n994 , n990 , n993 ); 
and ( n995 , n988 , n994 ); 
and ( n996 , n955 , n981 , n995 ); 
not ( n997 , n113 ); 
nor ( n998 , n996 , n997 ); 
nand ( n999 , n955 , n981 , n995 ); 
or ( n1000 , n999 , n113 ); 
nand ( n1001 , n1000 , n402 ); 
or ( n1002 , n998 , n1001 ); 
not ( n1003 , n114 ); 
or ( n1004 , n1003 , n402 ); 
nand ( n1005 , n1002 , n1004 ); 
not ( n1006 , n122 ); 
not ( n1007 , n1006 ); 
not ( n1008 , n788 ); 
not ( n1009 , n903 ); 
not ( n1010 , n847 ); 
nand ( n1011 , n1010 , n838 ); 
not ( n1012 , n882 ); 
or ( n1013 , n1011 , n1012 ); 
nor ( n1014 , n804 , n789 ); 
nand ( n1015 , n872 , n1014 ); 
nand ( n1016 , n1013 , n1015 ); 
not ( n1017 , n1016 ); 
or ( n1018 , n1009 , n1017 ); 
not ( n1019 , n906 ); 
not ( n1020 , n1014 ); 
nand ( n1021 , n1020 , n1011 ); 
nand ( n1022 , n1019 , n1021 , n778 ); 
nand ( n1023 , n1018 , n1022 ); 
nand ( n1024 , n1008 , n1023 ); 
nand ( n1025 , n963 , n915 ); 
and ( n1026 , n1024 , n887 , n949 , n1025 ); 
nand ( n1027 , n927 , n858 , n931 ); 
nand ( n1028 , n958 , n837 , n901 ); 
and ( n1029 , n1027 , n1028 ); 
and ( n1030 , n854 , n975 ); 
not ( n1031 , n872 ); 
nand ( n1032 , n810 , n1031 ); 
nor ( n1033 , n1032 , n880 ); 
nor ( n1034 , n1033 , n869 ); 
not ( n1035 , n1034 ); 
nand ( n1036 , n962 , n974 ); 
nand ( n1037 , n1036 , n831 ); 
nor ( n1038 , n1035 , n1037 ); 
nand ( n1039 , n1026 , n1029 , n1030 , n1038 ); 
not ( n1040 , n889 ); 
nor ( n1041 , n929 , n837 ); 
nand ( n1042 , n1040 , n1041 ); 
not ( n1043 , n1042 ); 
nor ( n1044 , n811 , n935 ); 
nand ( n1045 , n969 , n1044 ); 
not ( n1046 , n1045 ); 
nor ( n1047 , n1043 , n1046 ); 
nor ( n1048 , n978 , n993 ); 
nand ( n1049 , n1047 , n1048 ); 
not ( n1050 , n912 ); 
not ( n1051 , n1044 ); 
or ( n1052 , n1050 , n1051 ); 
nand ( n1053 , n1052 , n862 ); 
not ( n1054 , n1053 ); 
nand ( n1055 , n931 , n923 , n840 ); 
nand ( n1056 , n928 , n1055 ); 
not ( n1057 , n1056 ); 
nand ( n1058 , n1054 , n1057 ); 
nor ( n1059 , n1049 , n1058 ); 
nand ( n1060 , n1041 , n846 ); 
not ( n1061 , n1060 ); 
nand ( n1062 , n923 , n867 ); 
nor ( n1063 , n834 , n1062 ); 
nor ( n1064 , n1061 , n1063 ); 
nand ( n1065 , n1064 , n973 , n988 ); 
or ( n1066 , n912 , n1062 ); 
nand ( n1067 , n1066 , n943 ); 
not ( n1068 , n1067 ); 
nand ( n1069 , n920 , n1068 ); 
nor ( n1070 , n1065 , n1069 ); 
nand ( n1071 , n1059 , n1070 ); 
nor ( n1072 , n1039 , n1071 ); 
not ( n1073 , n1072 ); 
or ( n1074 , n1007 , n1073 ); 
nand ( n1075 , n1074 , n391 ); 
not ( n1076 , n1039 ); 
not ( n1077 , n1071 ); 
and ( n1078 , n1076 , n1077 ); 
nor ( n1079 , n1078 , n1006 ); 
or ( n1080 , n1075 , n1079 ); 
not ( n1081 , n123 ); 
or ( n1082 , n1081 , n391 ); 
nand ( n1083 , n1080 , n1082 ); 
and ( n1084 , n20 , n388 ); 
and ( n1085 , n3 , n21 ); 
nor ( n1086 , n1084 , n1085 ); 
and ( n1087 , n391 , n1086 ); 
not ( n1088 , n391 ); 
xor ( n1089 , n27 , n28 ); 
buf ( n1090 , n1089 ); 
not ( n1091 , n23 ); 
not ( n1092 , n24 ); 
not ( n1093 , n1092 ); 
or ( n1094 , n1091 , n1093 ); 
not ( n1095 , n23 ); 
nand ( n1096 , n24 , n1095 ); 
nand ( n1097 , n1094 , n1096 ); 
buf ( n1098 , n1097 ); 
not ( n1099 , n1098 ); 
not ( n1100 , n25 ); 
not ( n1101 , n26 ); 
not ( n1102 , n1101 ); 
or ( n1103 , n1100 , n1102 ); 
not ( n1104 , n25 ); 
nand ( n1105 , n1104 , n26 ); 
nand ( n1106 , n1103 , n1105 ); 
nand ( n1107 , n1099 , n1106 ); 
not ( n1108 , n1107 ); 
nand ( n1109 , n1090 , n1108 ); 
not ( n1110 , n1109 ); 
xor ( n1111 , n31 , n32 ); 
buf ( n1112 , n1111 ); 
and ( n1113 , n29 , n30 ); 
not ( n1114 , n29 ); 
not ( n1115 , n30 ); 
and ( n1116 , n1114 , n1115 ); 
nor ( n1117 , n1113 , n1116 ); 
not ( n1118 , n1117 ); 
buf ( n1119 , n1118 ); 
and ( n1120 , n33 , n34 ); 
not ( n1121 , n33 ); 
not ( n1122 , n34 ); 
and ( n1123 , n1121 , n1122 ); 
or ( n1124 , n1120 , n1123 ); 
not ( n1125 , n1124 ); 
nand ( n1126 , n1110 , n1112 , n1119 , n1125 ); 
not ( n1127 , n1126 ); 
not ( n1128 , n1124 ); 
buf ( n1129 , n1128 ); 
not ( n1130 , n1129 ); 
nor ( n1131 , n1098 , n1106 ); 
buf ( n1132 , n1131 ); 
not ( n1133 , n1089 ); 
nand ( n1134 , n1132 , n1133 , n1118 ); 
not ( n1135 , n1111 ); 
nor ( n1136 , n1134 , n1135 ); 
not ( n1137 , n1136 ); 
or ( n1138 , n1130 , n1137 ); 
not ( n1139 , n1128 ); 
not ( n1140 , n1111 ); 
not ( n1141 , n1140 ); 
nor ( n1142 , n1109 , n1119 ); 
nand ( n1143 , n1139 , n1141 , n1142 ); 
nand ( n1144 , n1138 , n1143 ); 
nor ( n1145 , n1127 , n1144 ); 
not ( n1146 , n1124 ); 
not ( n1147 , n1146 ); 
not ( n1148 , n1147 ); 
and ( n1149 , n1089 , n1131 ); 
buf ( n1150 , n1117 ); 
not ( n1151 , n1150 ); 
nand ( n1152 , n1149 , n1151 ); 
not ( n1153 , n1111 ); 
not ( n1154 , n1153 ); 
not ( n1155 , n1154 ); 
nor ( n1156 , n1152 , n1155 ); 
nand ( n1157 , n1148 , n1156 ); 
not ( n1158 , n1132 ); 
not ( n1159 , n1158 ); 
not ( n1160 , n1111 ); 
not ( n1161 , n1160 ); 
buf ( n1162 , n1117 ); 
buf ( n1163 , n1133 ); 
nand ( n1164 , n1159 , n1161 , n1162 , n1163 ); 
not ( n1165 , n1164 ); 
nand ( n1166 , n1165 , n1129 ); 
not ( n1167 , n1166 ); 
not ( n1168 , n1149 ); 
not ( n1169 , n1162 ); 
nor ( n1170 , n1168 , n1169 ); 
not ( n1171 , n1140 ); 
nand ( n1172 , n1170 , n1171 , n1146 ); 
not ( n1173 , n1172 ); 
nor ( n1174 , n1167 , n1173 ); 
buf ( n1175 , n1124 ); 
not ( n1176 , n1175 ); 
not ( n1177 , n1098 ); 
not ( n1178 , n1177 ); 
not ( n1179 , n1106 ); 
nand ( n1180 , n1178 , n1089 , n1150 , n1179 ); 
nor ( n1181 , n1154 , n1180 ); 
nand ( n1182 , n1176 , n1181 ); 
not ( n1183 , n1182 ); 
nor ( n1184 , n1164 , n1129 ); 
nor ( n1185 , n1183 , n1184 ); 
nand ( n1186 , n1145 , n1157 , n1174 , n1185 ); 
not ( n1187 , n1186 ); 
not ( n1188 , n1139 ); 
not ( n1189 , n1135 ); 
nand ( n1190 , n1132 , n1133 , n1162 ); 
nor ( n1191 , n1189 , n1190 ); 
and ( n1192 , n1188 , n1191 ); 
not ( n1193 , n1188 ); 
not ( n1194 , n1171 ); 
not ( n1195 , n1106 ); 
not ( n1196 , n1195 ); 
not ( n1197 , n1089 ); 
and ( n1198 , n29 , n30 ); 
not ( n1199 , n29 ); 
and ( n1200 , n1199 , n1115 ); 
nor ( n1201 , n1198 , n1200 ); 
nand ( n1202 , n1098 , n1201 ); 
or ( n1203 , n1196 , n1197 , n1202 ); 
buf ( n1204 , n1195 ); 
nor ( n1205 , n1098 , n1201 ); 
nand ( n1206 , n1197 , n1205 ); 
or ( n1207 , n1204 , n1206 ); 
nand ( n1208 , n1203 , n1207 ); 
not ( n1209 , n1208 ); 
or ( n1210 , n1194 , n1209 ); 
not ( n1211 , n1204 ); 
not ( n1212 , n1163 ); 
not ( n1213 , n1205 ); 
nand ( n1214 , n1213 , n1202 ); 
nand ( n1215 , n1211 , n1212 , n1135 , n1214 ); 
nand ( n1216 , n1210 , n1215 ); 
and ( n1217 , n1193 , n1216 ); 
nor ( n1218 , n1192 , n1217 ); 
not ( n1219 , n1153 ); 
not ( n1220 , n1219 ); 
not ( n1221 , n1195 ); 
and ( n1222 , n1150 , n1197 , n1221 , n1177 ); 
nand ( n1223 , n1220 , n1222 ); 
not ( n1224 , n1223 ); 
nand ( n1225 , n1148 , n1224 ); 
nand ( n1226 , n1170 , n1155 , n1175 ); 
and ( n1227 , n1132 , n1151 , n1133 , n1153 ); 
nand ( n1228 , n1148 , n1227 ); 
nand ( n1229 , n1218 , n1225 , n1226 , n1228 ); 
nand ( n1230 , n1098 , n1106 ); 
nor ( n1231 , n1150 , n1197 , n1230 ); 
nand ( n1232 , n1155 , n1231 ); 
nor ( n1233 , n1130 , n1232 ); 
not ( n1234 , n1125 ); 
not ( n1235 , n1234 ); 
nor ( n1236 , n1152 , n1112 ); 
not ( n1237 , n1236 ); 
or ( n1238 , n1235 , n1237 ); 
nor ( n1239 , n1230 , n1089 ); 
and ( n1240 , n1162 , n1239 ); 
nand ( n1241 , n1240 , n1220 , n1125 ); 
nand ( n1242 , n1238 , n1241 ); 
nor ( n1243 , n1233 , n1242 ); 
not ( n1244 , n1089 ); 
nand ( n1245 , n1195 , n1098 , n1244 ); 
not ( n1246 , n1245 ); 
nand ( n1247 , n1162 , n1246 ); 
nor ( n1248 , n1247 , n1112 ); 
nand ( n1249 , n1148 , n1248 ); 
nand ( n1250 , n1142 , n1220 , n1176 ); 
nand ( n1251 , n1239 , n1151 ); 
nor ( n1252 , n1251 , n1219 ); 
nand ( n1253 , n1175 , n1252 ); 
nand ( n1254 , n1250 , n1253 ); 
nand ( n1255 , n1181 , n1234 ); 
not ( n1256 , n1201 ); 
nand ( n1257 , n1178 , n1089 , n1256 , n1179 ); 
nor ( n1258 , n1219 , n1257 ); 
nand ( n1259 , n1234 , n1258 ); 
nand ( n1260 , n1255 , n1259 ); 
nor ( n1261 , n1254 , n1260 ); 
nand ( n1262 , n1243 , n1249 , n1261 ); 
nor ( n1263 , n1229 , n1262 ); 
not ( n1264 , n1230 ); 
nand ( n1265 , n1264 , n1162 , n1111 , n1090 ); 
not ( n1266 , n1265 ); 
nand ( n1267 , n1129 , n1266 ); 
not ( n1268 , n1257 ); 
nand ( n1269 , n1141 , n1268 ); 
not ( n1270 , n1269 ); 
not ( n1271 , n1135 ); 
not ( n1272 , n1251 ); 
nand ( n1273 , n1271 , n1272 ); 
not ( n1274 , n1273 ); 
or ( n1275 , n1270 , n1274 ); 
nand ( n1276 , n1275 , n1188 ); 
nand ( n1277 , n1267 , n1276 ); 
nand ( n1278 , n1161 , n1169 , n1246 ); 
nor ( n1279 , n1175 , n1278 ); 
not ( n1280 , n1279 ); 
not ( n1281 , n1139 ); 
nor ( n1282 , n1281 , n1223 ); 
not ( n1283 , n1282 ); 
nand ( n1284 , n1280 , n1283 ); 
not ( n1285 , n1139 ); 
nor ( n1286 , n1285 , n1265 ); 
not ( n1287 , n1286 ); 
not ( n1288 , n1140 ); 
nand ( n1289 , n1175 , n1288 , n1240 ); 
nor ( n1290 , n1125 , n1278 ); 
not ( n1291 , n1290 ); 
nand ( n1292 , n1287 , n1289 , n1291 ); 
nor ( n1293 , n1277 , n1284 , n1292 ); 
nand ( n1294 , n1187 , n1263 , n1293 ); 
not ( n1295 , n22 ); 
and ( n1296 , n1294 , n1295 ); 
not ( n1297 , n1294 ); 
and ( n1298 , n1297 , n22 ); 
nor ( n1299 , n1296 , n1298 ); 
and ( n1300 , n1088 , n1299 ); 
nor ( n1301 , n1087 , n1300 ); 
and ( n1302 , n35 , n388 ); 
and ( n1303 , n3 , n36 ); 
nor ( n1304 , n1302 , n1303 ); 
and ( n1305 , n402 , n1304 ); 
not ( n1306 , n402 ); 
not ( n1307 , n1180 ); 
nand ( n1308 , n1307 , n1288 , n1125 ); 
not ( n1309 , n1247 ); 
nand ( n1310 , n1129 , n1288 , n1309 ); 
and ( n1311 , n1276 , n1308 , n1310 ); 
and ( n1312 , n1176 , n1141 , n1231 ); 
nor ( n1313 , n1312 , n1286 ); 
nor ( n1314 , n1282 , n1290 ); 
nand ( n1315 , n1311 , n1313 , n1314 ); 
not ( n1316 , n1188 ); 
not ( n1317 , n1140 ); 
nand ( n1318 , n1317 , n1222 ); 
not ( n1319 , n1318 ); 
not ( n1320 , n1319 ); 
or ( n1321 , n1316 , n1320 ); 
nand ( n1322 , n1321 , n1166 ); 
nor ( n1323 , n1322 , n1144 ); 
not ( n1324 , n1127 ); 
nor ( n1325 , n1318 , n1129 ); 
not ( n1326 , n1325 ); 
nand ( n1327 , n1324 , n1326 ); 
not ( n1328 , n1182 ); 
not ( n1329 , n1328 ); 
nand ( n1330 , n1156 , n1147 ); 
nand ( n1331 , n1329 , n1330 ); 
nor ( n1332 , n1327 , n1331 ); 
nand ( n1333 , n1323 , n1332 ); 
nor ( n1334 , n1315 , n1333 ); 
and ( n1335 , n1129 , n1236 ); 
not ( n1336 , n1129 ); 
and ( n1337 , n1336 , n1227 ); 
nor ( n1338 , n1335 , n1337 ); 
not ( n1339 , n1338 ); 
nor ( n1340 , n1339 , n1233 ); 
not ( n1341 , n1250 ); 
nand ( n1342 , n1119 , n1246 ); 
nor ( n1343 , n1342 , n1171 , n1175 ); 
not ( n1344 , n1343 ); 
nand ( n1345 , n1175 , n1248 ); 
nand ( n1346 , n1344 , n1345 ); 
nor ( n1347 , n1341 , n1346 ); 
not ( n1348 , n1252 ); 
nor ( n1349 , n1348 , n1130 ); 
nand ( n1350 , n1253 , n1259 ); 
nor ( n1351 , n1349 , n1350 ); 
nand ( n1352 , n1340 , n1347 , n1351 ); 
not ( n1353 , n1139 ); 
nor ( n1354 , n1090 , n1107 ); 
nand ( n1355 , n1169 , n1354 ); 
nor ( n1356 , n1141 , n1355 ); 
and ( n1357 , n1353 , n1356 ); 
not ( n1358 , n1353 ); 
nand ( n1359 , n1230 , n1158 ); 
nand ( n1360 , n1359 , n1163 , n1135 , n1162 ); 
or ( n1361 , n1118 , n1132 ); 
nor ( n1362 , n1133 , n1160 ); 
nand ( n1363 , n1118 , n1230 ); 
nand ( n1364 , n1361 , n1362 , n1363 ); 
nand ( n1365 , n1360 , n1364 ); 
and ( n1366 , n1358 , n1365 ); 
nor ( n1367 , n1357 , n1366 ); 
nand ( n1368 , n1367 , n1226 , n1228 ); 
nor ( n1369 , n1352 , n1368 ); 
nand ( n1370 , n1334 , n1369 ); 
not ( n1371 , n37 ); 
and ( n1372 , n1370 , n1371 ); 
not ( n1373 , n1370 ); 
and ( n1374 , n1373 , n37 ); 
nor ( n1375 , n1372 , n1374 ); 
and ( n1376 , n1306 , n1375 ); 
nor ( n1377 , n1305 , n1376 ); 
and ( n1378 , n56 , n388 ); 
and ( n1379 , n3 , n57 ); 
nor ( n1380 , n1378 , n1379 ); 
and ( n1381 , n402 , n1380 ); 
not ( n1382 , n402 ); 
not ( n1383 , n13 ); 
and ( n1384 , n14 , n1383 ); 
not ( n1385 , n14 ); 
and ( n1386 , n1385 , n13 ); 
nor ( n1387 , n1384 , n1386 ); 
buf ( n1388 , n1387 ); 
buf ( n1389 , n1388 ); 
not ( n1390 , n15 ); 
and ( n1391 , n16 , n1390 ); 
not ( n1392 , n16 ); 
and ( n1393 , n1392 , n15 ); 
nor ( n1394 , n1391 , n1393 ); 
not ( n1395 , n1394 ); 
not ( n1396 , n1395 ); 
not ( n1397 , n1396 ); 
and ( n1398 , n6 , n5 ); 
not ( n1399 , n6 ); 
not ( n1400 , n5 ); 
and ( n1401 , n1399 , n1400 ); 
nor ( n1402 , n1398 , n1401 ); 
not ( n1403 , n1402 ); 
not ( n1404 , n1403 ); 
xor ( n1405 , n9 , n10 ); 
and ( n1406 , n8 , n7 ); 
not ( n1407 , n8 ); 
not ( n1408 , n7 ); 
and ( n1409 , n1407 , n1408 ); 
nor ( n1410 , n1406 , n1409 ); 
not ( n1411 , n1410 ); 
nand ( n1412 , n1404 , n1405 , n1411 ); 
not ( n1413 , n11 ); 
not ( n1414 , n12 ); 
not ( n1415 , n1414 ); 
or ( n1416 , n1413 , n1415 ); 
not ( n1417 , n11 ); 
nand ( n1418 , n12 , n1417 ); 
nand ( n1419 , n1416 , n1418 ); 
buf ( n1420 , n1419 ); 
buf ( n1421 , n1420 ); 
nor ( n1422 , n1412 , n1421 ); 
nand ( n1423 , n1389 , n1397 , n1422 ); 
buf ( n1424 , n1394 ); 
buf ( n1425 , n1424 ); 
nor ( n1426 , n1410 , n1402 ); 
not ( n1427 , n1426 ); 
xnor ( n1428 , n10 , n9 ); 
not ( n1429 , n1428 ); 
not ( n1430 , n1429 ); 
nor ( n1431 , n1427 , n1430 ); 
buf ( n1432 , n1420 ); 
not ( n1433 , n1432 ); 
nand ( n1434 , n1431 , n1388 , n1433 ); 
nor ( n1435 , n1425 , n1434 ); 
not ( n1436 , n1435 ); 
and ( n1437 , n1423 , n1436 ); 
buf ( n1438 , n1424 ); 
nand ( n1439 , n1420 , n1387 ); 
nor ( n1440 , n1439 , n1412 ); 
nand ( n1441 , n1438 , n1440 ); 
buf ( n1442 , n1420 ); 
not ( n1443 , n1442 ); 
not ( n1444 , n1403 ); 
not ( n1445 , n1444 ); 
nand ( n1446 , n1445 , n1405 , n1410 ); 
nor ( n1447 , n1443 , n1446 ); 
not ( n1448 , n1388 ); 
not ( n1449 , n1448 ); 
nand ( n1450 , n1447 , n1449 , n1425 ); 
buf ( n1451 , n1394 ); 
not ( n1452 , n1451 ); 
buf ( n1453 , n1420 ); 
buf ( n1454 , n1402 ); 
not ( n1455 , n1454 ); 
buf ( n1456 , n1410 ); 
nand ( n1457 , n1455 , n1456 , n1428 ); 
nor ( n1458 , n1453 , n1457 ); 
nand ( n1459 , n1389 , n1452 , n1458 ); 
and ( n1460 , n1441 , n1450 , n1459 ); 
not ( n1461 , n1446 ); 
not ( n1462 , n1421 ); 
nand ( n1463 , n1461 , n1397 , n1449 , n1462 ); 
not ( n1464 , n1463 ); 
not ( n1465 , n1464 ); 
not ( n1466 , n1387 ); 
not ( n1467 , n1466 ); 
nand ( n1468 , n1454 , n1410 ); 
nor ( n1469 , n1468 , n1405 ); 
nand ( n1470 , n1467 , n1451 , n1443 , n1469 ); 
and ( n1471 , n1428 , n1454 , n1411 ); 
not ( n1472 , n1471 ); 
not ( n1473 , n1472 ); 
not ( n1474 , n13 ); 
not ( n1475 , n14 ); 
not ( n1476 , n1475 ); 
or ( n1477 , n1474 , n1476 ); 
nand ( n1478 , n14 , n1383 ); 
nand ( n1479 , n1477 , n1478 ); 
nor ( n1480 , n1420 , n1479 ); 
nand ( n1481 , n1473 , n1480 , n1396 ); 
and ( n1482 , n1470 , n1481 ); 
nand ( n1483 , n1437 , n1460 , n1465 , n1482 ); 
not ( n1484 , n1394 ); 
nor ( n1485 , n1484 , n1479 ); 
nand ( n1486 , n1485 , n1453 , n1431 ); 
not ( n1487 , n1486 ); 
not ( n1488 , n1403 ); 
not ( n1489 , n1488 ); 
nor ( n1490 , n1489 , n1484 ); 
not ( n1491 , n1490 ); 
not ( n1492 , n1404 ); 
nand ( n1493 , n1492 , n1484 ); 
nand ( n1494 , n1491 , n1493 ); 
not ( n1495 , n1429 ); 
nand ( n1496 , n1494 , n1495 , n1388 ); 
not ( n1497 , n1456 ); 
not ( n1498 , n1497 ); 
not ( n1499 , n1498 ); 
not ( n1500 , n1432 ); 
not ( n1501 , n1500 ); 
not ( n1502 , n1501 ); 
nor ( n1503 , n1496 , n1499 , n1502 ); 
nor ( n1504 , n1487 , n1503 ); 
not ( n1505 , n1425 ); 
buf ( n1506 , n1479 ); 
not ( n1507 , n1420 ); 
not ( n1508 , n1507 ); 
nand ( n1509 , n1454 , n1405 , n1410 ); 
not ( n1510 , n1509 ); 
and ( n1511 , n1506 , n1508 , n1510 ); 
nand ( n1512 , n1505 , n1511 ); 
not ( n1513 , n1512 ); 
not ( n1514 , n1424 ); 
buf ( n1515 , n1514 ); 
not ( n1516 , n1420 ); 
nand ( n1517 , n1428 , n1426 ); 
nor ( n1518 , n1516 , n1517 ); 
nand ( n1519 , n1389 , n1518 ); 
nor ( n1520 , n1515 , n1519 ); 
nor ( n1521 , n1513 , n1520 ); 
not ( n1522 , n1514 ); 
not ( n1523 , n1421 ); 
not ( n1524 , n1446 ); 
nand ( n1525 , n1523 , n1524 ); 
not ( n1526 , n1479 ); 
not ( n1527 , n1526 ); 
buf ( n1528 , n1527 ); 
nor ( n1529 , n1525 , n1528 ); 
nand ( n1530 , n1522 , n1529 ); 
not ( n1531 , n1489 ); 
or ( n1532 , n1531 , n1495 , n1395 ); 
nand ( n1533 , n1404 , n1428 ); 
or ( n1534 , n1396 , n1533 ); 
nand ( n1535 , n1532 , n1534 ); 
nand ( n1536 , n1528 , n1499 , n1502 , n1535 ); 
nand ( n1537 , n1504 , n1521 , n1530 , n1536 ); 
nor ( n1538 , n1483 , n1537 ); 
not ( n1539 , n1396 ); 
not ( n1540 , n1526 ); 
and ( n1541 , n1469 , n1421 , n1540 ); 
nand ( n1542 , n1539 , n1541 ); 
not ( n1543 , n1422 ); 
nor ( n1544 , n1389 , n1543 ); 
nand ( n1545 , n1539 , n1544 ); 
nand ( n1546 , n1542 , n1545 ); 
nand ( n1547 , n1528 , n1397 , n1447 ); 
not ( n1548 , n1427 ); 
not ( n1549 , n1526 ); 
nand ( n1550 , n1548 , n1549 , n1442 , n1405 ); 
not ( n1551 , n1550 ); 
nand ( n1552 , n1539 , n1551 ); 
nand ( n1553 , n1547 , n1552 ); 
nor ( n1554 , n1546 , n1553 ); 
buf ( n1555 , n1451 ); 
nand ( n1556 , n1555 , n1511 ); 
not ( n1557 , n1556 ); 
buf ( n1558 , n1420 ); 
nand ( n1559 , n1558 , n1471 ); 
not ( n1560 , n1559 ); 
nand ( n1561 , n1528 , n1560 ); 
nor ( n1562 , n1515 , n1561 ); 
nor ( n1563 , n1557 , n1562 ); 
not ( n1564 , n1412 ); 
nand ( n1565 , n1564 , n1425 , n1528 , n1500 ); 
not ( n1566 , n1565 ); 
and ( n1567 , n1469 , n1516 , n1506 ); 
nand ( n1568 , n1539 , n1567 ); 
not ( n1569 , n1568 ); 
nor ( n1570 , n1566 , n1569 ); 
nand ( n1571 , n1554 , n1563 , n1570 ); 
buf ( n1572 , n1506 ); 
not ( n1573 , n1424 ); 
nand ( n1574 , n1572 , n1573 , n1518 ); 
not ( n1575 , n1574 ); 
nor ( n1576 , n1517 , n1442 ); 
not ( n1577 , n1526 ); 
and ( n1578 , n1576 , n1577 , n1451 ); 
nor ( n1579 , n1575 , n1578 ); 
nand ( n1580 , n1505 , n1440 ); 
not ( n1581 , n1442 ); 
and ( n1582 , n1524 , n1581 , n1577 ); 
nand ( n1583 , n1505 , n1582 ); 
and ( n1584 , n1579 , n1580 , n1583 ); 
not ( n1585 , n1539 ); 
nor ( n1586 , n1572 , n1559 ); 
not ( n1587 , n1586 ); 
or ( n1588 , n1585 , n1587 ); 
and ( n1589 , n1388 , n1433 , n1510 ); 
nand ( n1590 , n1539 , n1589 ); 
nand ( n1591 , n1588 , n1590 ); 
not ( n1592 , n1591 ); 
not ( n1593 , n1457 ); 
buf ( n1594 , n1420 ); 
nand ( n1595 , n1593 , n1528 , n1438 , n1594 ); 
not ( n1596 , n1595 ); 
and ( n1597 , n1528 , n1555 , n1458 ); 
nor ( n1598 , n1596 , n1597 ); 
nand ( n1599 , n1584 , n1592 , n1598 ); 
nor ( n1600 , n1571 , n1599 ); 
nand ( n1601 , n1538 , n1600 ); 
not ( n1602 , n58 ); 
and ( n1603 , n1601 , n1602 ); 
not ( n1604 , n1601 ); 
and ( n1605 , n1604 , n58 ); 
nor ( n1606 , n1603 , n1605 ); 
and ( n1607 , n1382 , n1606 ); 
nor ( n1608 , n1381 , n1607 ); 
nand ( n1609 , n290 , n268 ); 
not ( n1610 , n1609 ); 
nor ( n1611 , n377 , n1610 ); 
not ( n1612 , n317 ); 
nand ( n1613 , n1612 , n362 ); 
not ( n1614 , n292 ); 
and ( n1615 , n1611 , n1613 , n1614 , n303 ); 
not ( n1616 , n178 ); 
nand ( n1617 , n1616 , n212 ); 
and ( n1618 , n1617 , n270 ); 
not ( n1619 , n260 ); 
not ( n1620 , n264 ); 
or ( n1621 , n1619 , n1620 ); 
nand ( n1622 , n1621 , n223 ); 
not ( n1623 , n1622 ); 
nor ( n1624 , n225 , n243 ); 
not ( n1625 , n1624 ); 
nand ( n1626 , n1618 , n1623 , n234 , n1625 ); 
nand ( n1627 , n257 , n332 ); 
nor ( n1628 , n1626 , n1627 ); 
nand ( n1629 , n1615 , n1628 ); 
not ( n1630 , n1629 ); 
nor ( n1631 , n241 , n230 ); 
nand ( n1632 , n277 , n238 , n1631 ); 
nand ( n1633 , n201 , n214 ); 
not ( n1634 , n1633 ); 
nand ( n1635 , n182 , n1634 ); 
not ( n1636 , n189 ); 
nor ( n1637 , n1636 , n201 ); 
nand ( n1638 , n250 , n1637 ); 
nand ( n1639 , n1635 , n1638 ); 
not ( n1640 , n341 ); 
nor ( n1641 , n259 , n1640 ); 
nand ( n1642 , n1639 , n211 , n1641 ); 
nand ( n1643 , n1632 , n1642 ); 
not ( n1644 , n1643 ); 
not ( n1645 , n320 ); 
nand ( n1646 , n296 , n307 ); 
not ( n1647 , n1646 ); 
and ( n1648 , n1645 , n1647 ); 
not ( n1649 , n216 ); 
not ( n1650 , n307 ); 
nand ( n1651 , n1649 , n1650 ); 
not ( n1652 , n1651 ); 
and ( n1653 , n1652 , n230 ); 
nor ( n1654 , n1648 , n1653 ); 
not ( n1655 , n1640 ); 
nand ( n1656 , n327 , n178 ); 
nor ( n1657 , n1654 , n1655 , n1656 ); 
nor ( n1658 , n370 , n1657 ); 
nand ( n1659 , n290 , n310 ); 
nand ( n1660 , n301 , n236 ); 
nand ( n1661 , n1644 , n1658 , n1659 , n1660 ); 
nand ( n1662 , n277 , n379 ); 
not ( n1663 , n1662 ); 
nor ( n1664 , n1616 , n316 ); 
nor ( n1665 , n1663 , n1664 ); 
nand ( n1666 , n365 , n248 , n277 ); 
and ( n1667 , n1666 , n328 ); 
not ( n1668 , n178 ); 
nand ( n1669 , n1668 , n375 ); 
and ( n1670 , n1669 , n330 ); 
nor ( n1671 , n225 , n322 ); 
nor ( n1672 , n312 , n1671 ); 
nand ( n1673 , n1665 , n1667 , n1670 , n1672 ); 
nor ( n1674 , n1661 , n1673 ); 
and ( n1675 , n1630 , n282 , n1674 ); 
not ( n1676 , n60 ); 
nor ( n1677 , n1675 , n1676 ); 
not ( n1678 , n1676 ); 
nand ( n1679 , n282 , n1674 ); 
nor ( n1680 , n1629 , n1679 ); 
not ( n1681 , n1680 ); 
or ( n1682 , n1678 , n1681 ); 
not ( n1683 , n391 ); 
nand ( n1684 , n1682 , n1683 ); 
or ( n1685 , n1677 , n1684 ); 
and ( n1686 , n59 , n388 ); 
and ( n1687 , n3 , n38 ); 
nor ( n1688 , n1686 , n1687 ); 
or ( n1689 , n1688 , n631 ); 
nand ( n1690 , n1685 , n1689 ); 
not ( n1691 , n402 ); 
not ( n1692 , n74 ); 
and ( n1693 , n1691 , n1692 ); 
not ( n1694 , n1691 ); 
and ( n1695 , n1694 , n1299 ); 
nor ( n1696 , n1693 , n1695 ); 
not ( n1697 , n776 ); 
not ( n1698 , n805 ); 
and ( n1699 , n1697 , n1698 ); 
and ( n1700 , n872 , n924 ); 
nor ( n1701 , n1699 , n1700 ); 
not ( n1702 , n809 ); 
nand ( n1703 , n1702 , n838 ); 
or ( n1704 , n1701 , n1703 ); 
or ( n1705 , n906 , n1015 ); 
nand ( n1706 , n1704 , n1705 ); 
nand ( n1707 , n788 , n1706 ); 
nand ( n1708 , n937 , n822 , n1707 ); 
not ( n1709 , n899 ); 
nand ( n1710 , n850 , n833 , n951 , n1709 ); 
nand ( n1711 , n1710 , n1027 , n932 ); 
nor ( n1712 , n1708 , n1711 ); 
nor ( n1713 , n993 , n855 ); 
and ( n1714 , n1040 , n853 ); 
not ( n1715 , n1028 ); 
nor ( n1716 , n1714 , n1715 ); 
nand ( n1717 , n1716 , n813 , n1034 ); 
not ( n1718 , n1717 ); 
and ( n1719 , n1712 , n1713 , n1718 ); 
not ( n1720 , n920 ); 
nor ( n1721 , n1720 , n1067 ); 
and ( n1722 , n970 , n967 ); 
not ( n1723 , n970 ); 
and ( n1724 , n1723 , n915 ); 
nor ( n1725 , n1722 , n1724 ); 
nand ( n1726 , n895 , n986 ); 
nor ( n1727 , n971 , n1726 ); 
nand ( n1728 , n1721 , n1725 , n1727 ); 
not ( n1729 , n1055 ); 
not ( n1730 , n834 ); 
not ( n1731 , n991 ); 
or ( n1732 , n1730 , n1731 ); 
nand ( n1733 , n1732 , n952 ); 
nor ( n1734 , n1729 , n1733 ); 
not ( n1735 , n983 ); 
nor ( n1736 , n964 , n1735 ); 
nand ( n1737 , n1040 , n985 ); 
nand ( n1738 , n1042 , n1045 , n1737 ); 
not ( n1739 , n1738 ); 
nand ( n1740 , n1734 , n1736 , n1739 ); 
nor ( n1741 , n1728 , n1740 ); 
nand ( n1742 , n1719 , n1741 ); 
or ( n1743 , n97 , n1742 ); 
nand ( n1744 , n1743 , n402 ); 
and ( n1745 , n1719 , n1741 ); 
not ( n1746 , n97 ); 
nor ( n1747 , n1745 , n1746 ); 
or ( n1748 , n1744 , n1747 ); 
not ( n1749 , n106 ); 
or ( n1750 , n1749 , n402 ); 
nand ( n1751 , n1748 , n1750 ); 
not ( n1752 , n135 ); 
not ( n1753 , n1752 ); 
not ( n1754 , n1148 ); 
not ( n1755 , n1754 ); 
not ( n1756 , n1212 ); 
not ( n1757 , n1756 ); 
and ( n1758 , n1196 , n1160 , n1205 ); 
not ( n1759 , n1758 ); 
nand ( n1760 , n1204 , n1154 , n1214 ); 
nand ( n1761 , n1759 , n1760 ); 
not ( n1762 , n1761 ); 
or ( n1763 , n1757 , n1762 ); 
nand ( n1764 , n1763 , n1232 ); 
not ( n1765 , n1764 ); 
or ( n1766 , n1755 , n1765 ); 
nand ( n1767 , n1766 , n1267 ); 
not ( n1768 , n1308 ); 
not ( n1769 , n1768 ); 
nand ( n1770 , n1769 , n1283 ); 
nor ( n1771 , n1767 , n1770 ); 
not ( n1772 , n1288 ); 
and ( n1773 , n1119 , n1110 ); 
nand ( n1774 , n1188 , n1772 , n1773 ); 
nand ( n1775 , n1250 , n1774 , n1338 ); 
nand ( n1776 , n1129 , n1191 ); 
not ( n1777 , n1776 ); 
not ( n1778 , n1345 ); 
nor ( n1779 , n1777 , n1778 ); 
not ( n1780 , n1350 ); 
nand ( n1781 , n1779 , n1255 , n1780 ); 
nor ( n1782 , n1775 , n1781 ); 
nand ( n1783 , n1771 , n1782 ); 
not ( n1784 , n1146 ); 
nor ( n1785 , n1355 , n1140 ); 
not ( n1786 , n1785 ); 
or ( n1787 , n1784 , n1786 ); 
nand ( n1788 , n1787 , n1126 ); 
nor ( n1789 , n1286 , n1788 ); 
not ( n1790 , n1273 ); 
nand ( n1791 , n1790 , n1147 ); 
nor ( n1792 , n1312 , n1279 ); 
not ( n1793 , n1172 ); 
nor ( n1794 , n1793 , n1290 ); 
and ( n1795 , n1789 , n1791 , n1792 , n1794 ); 
not ( n1796 , n1258 ); 
nor ( n1797 , n1147 , n1796 ); 
nor ( n1798 , n1349 , n1797 ); 
not ( n1799 , n1242 ); 
nand ( n1800 , n1798 , n1799 ); 
nand ( n1801 , n1129 , n1136 ); 
not ( n1802 , n1801 ); 
nor ( n1803 , n1802 , n1325 ); 
not ( n1804 , n1184 ); 
nand ( n1805 , n1803 , n1330 , n1804 ); 
nor ( n1806 , n1800 , n1805 ); 
nand ( n1807 , n1795 , n1806 ); 
nor ( n1808 , n1783 , n1807 ); 
not ( n1809 , n1808 ); 
or ( n1810 , n1753 , n1809 ); 
nand ( n1811 , n1810 , n402 ); 
not ( n1812 , n1807 ); 
and ( n1813 , n1812 , n1771 , n1782 ); 
nor ( n1814 , n1813 , n1752 ); 
or ( n1815 , n1811 , n1814 ); 
not ( n1816 , n136 ); 
or ( n1817 , n1816 , n402 ); 
nand ( n1818 , n1815 , n1817 ); 
not ( n1819 , n110 ); 
and ( n1820 , n1691 , n1819 ); 
not ( n1821 , n1691 ); 
and ( n1822 , n1821 , n1375 ); 
nor ( n1823 , n1820 , n1822 ); 
not ( n1824 , n368 ); 
not ( n1825 , n281 ); 
nor ( n1826 , n1824 , n1825 ); 
and ( n1827 , n380 , n1609 ); 
nand ( n1828 , n1826 , n1613 , n1827 ); 
not ( n1829 , n1828 ); 
not ( n1830 , n317 ); 
and ( n1831 , n320 , n1646 ); 
not ( n1832 , n320 ); 
and ( n1833 , n1832 , n1651 ); 
nor ( n1834 , n1831 , n1833 ); 
and ( n1835 , n1834 , n248 , n1655 ); 
not ( n1836 , n345 ); 
nand ( n1837 , n1836 , n342 ); 
nand ( n1838 , n1837 , n237 ); 
not ( n1839 , n356 ); 
nor ( n1840 , n1838 , n1839 , n336 ); 
nor ( n1841 , n1835 , n1840 ); 
or ( n1842 , n1830 , n1841 ); 
nand ( n1843 , n1842 , n1617 , n232 ); 
not ( n1844 , n372 ); 
not ( n1845 , n1844 ); 
not ( n1846 , n263 ); 
nand ( n1847 , n1846 , n364 ); 
nand ( n1848 , n1845 , n1847 ); 
nor ( n1849 , n1843 , n1848 ); 
not ( n1850 , n1660 ); 
nand ( n1851 , n1616 , n211 , n331 ); 
nand ( n1852 , n276 , n1851 ); 
nor ( n1853 , n1850 , n1852 ); 
nand ( n1854 , n1829 , n1849 , n1853 ); 
not ( n1855 , n1854 ); 
not ( n1856 , n271 ); 
nor ( n1857 , n311 , n236 ); 
not ( n1858 , n1857 ); 
not ( n1859 , n213 ); 
nor ( n1860 , n1859 , n318 ); 
nand ( n1861 , n1856 , n1858 , n1860 ); 
nand ( n1862 , n1625 , n1667 ); 
nor ( n1863 , n1861 , n1862 ); 
nand ( n1864 , n246 , n211 , n1631 ); 
and ( n1865 , n330 , n1864 ); 
and ( n1866 , n1865 , n293 , n1665 , n315 ); 
nand ( n1867 , n1863 , n1866 ); 
not ( n1868 , n1867 ); 
and ( n1869 , n1855 , n1868 ); 
not ( n1870 , n118 ); 
nor ( n1871 , n1869 , n1870 ); 
not ( n1872 , n1870 ); 
nor ( n1873 , n1854 , n1867 ); 
not ( n1874 , n1873 ); 
or ( n1875 , n1872 , n1874 ); 
nand ( n1876 , n1875 , n402 ); 
or ( n1877 , n1871 , n1876 ); 
not ( n1878 , n119 ); 
or ( n1879 , n1878 , n402 ); 
nand ( n1880 , n1877 , n1879 ); 
not ( n1881 , n120 ); 
not ( n1882 , n1881 ); 
and ( n1883 , n16 , n95 ); 
not ( n1884 , n16 ); 
not ( n1885 , n95 ); 
and ( n1886 , n1884 , n1885 ); 
nor ( n1887 , n1883 , n1886 ); 
buf ( n1888 , n1887 ); 
not ( n1889 , n1888 ); 
not ( n1890 , n1889 ); 
not ( n1891 , n1890 ); 
xor ( n1892 , n14 , n94 ); 
not ( n1893 , n1892 ); 
not ( n1894 , n1893 ); 
not ( n1895 , n1894 ); 
not ( n1896 , n90 ); 
not ( n1897 , n91 ); 
not ( n1898 , n1897 ); 
or ( n1899 , n1896 , n1898 ); 
not ( n1900 , n90 ); 
nand ( n1901 , n91 , n1900 ); 
nand ( n1902 , n1899 , n1901 ); 
not ( n1903 , n1902 ); 
xor ( n1904 , n88 , n89 ); 
not ( n1905 , n92 ); 
not ( n1906 , n24 ); 
not ( n1907 , n1906 ); 
or ( n1908 , n1905 , n1907 ); 
not ( n1909 , n92 ); 
nand ( n1910 , n1909 , n24 ); 
nand ( n1911 , n1908 , n1910 ); 
buf ( n1912 , n1911 ); 
nand ( n1913 , n1903 , n1904 , n1912 ); 
xor ( n1914 , n26 , n93 ); 
buf ( n1915 , n1914 ); 
not ( n1916 , n1915 ); 
nor ( n1917 , n1913 , n1916 ); 
not ( n1918 , n1917 ); 
nor ( n1919 , n1895 , n1918 ); 
nand ( n1920 , n1891 , n1919 ); 
not ( n1921 , n1920 ); 
not ( n1922 , n1889 ); 
not ( n1923 , n1903 ); 
not ( n1924 , n1912 ); 
not ( n1925 , n1904 ); 
and ( n1926 , n1923 , n1924 , n1925 ); 
not ( n1927 , n1926 ); 
not ( n1928 , n1915 ); 
nor ( n1929 , n1927 , n1928 ); 
nand ( n1930 , n1929 , n1895 ); 
nor ( n1931 , n1922 , n1930 ); 
nor ( n1932 , n1921 , n1931 ); 
not ( n1933 , n1913 ); 
not ( n1934 , n1914 ); 
nor ( n1935 , n1892 , n1887 ); 
nand ( n1936 , n1934 , n1935 ); 
not ( n1937 , n1936 ); 
and ( n1938 , n1933 , n1937 ); 
buf ( n1939 , n1888 ); 
not ( n1940 , n1939 ); 
buf ( n1941 , n1893 ); 
not ( n1942 , n1941 ); 
not ( n1943 , n1914 ); 
not ( n1944 , n1943 ); 
not ( n1945 , n1902 ); 
xor ( n1946 , n88 , n89 ); 
nand ( n1947 , n1945 , n1946 ); 
nor ( n1948 , n1912 , n1947 ); 
nand ( n1949 , n1944 , n1948 ); 
nor ( n1950 , n1942 , n1949 ); 
nand ( n1951 , n1940 , n1950 ); 
not ( n1952 , n1951 ); 
nor ( n1953 , n1938 , n1952 ); 
not ( n1954 , n1939 ); 
buf ( n1955 , n1893 ); 
not ( n1956 , n1955 ); 
not ( n1957 , n1949 ); 
nand ( n1958 , n1954 , n1956 , n1957 ); 
not ( n1959 , n1958 ); 
buf ( n1960 , n1923 ); 
not ( n1961 , n1912 ); 
not ( n1962 , n1961 ); 
nand ( n1963 , n1904 , n1914 ); 
not ( n1964 , n1963 ); 
nand ( n1965 , n1962 , n1964 , n1935 ); 
not ( n1966 , n1904 ); 
not ( n1967 , n1966 ); 
not ( n1968 , n1934 ); 
or ( n1969 , n1967 , n1968 ); 
nand ( n1970 , n1969 , n1963 ); 
not ( n1971 , n1893 ); 
not ( n1972 , n1887 ); 
nor ( n1973 , n1912 , n1972 ); 
nand ( n1974 , n1970 , n1971 , n1973 ); 
nand ( n1975 , n1965 , n1974 ); 
and ( n1976 , n1960 , n1975 ); 
nor ( n1977 , n1959 , n1976 ); 
and ( n1978 , n1932 , n1953 , n1977 ); 
not ( n1979 , n1941 ); 
not ( n1980 , n1979 ); 
not ( n1981 , n1916 ); 
not ( n1982 , n1912 ); 
nand ( n1983 , n1946 , n1902 ); 
nor ( n1984 , n1982 , n1983 ); 
nand ( n1985 , n1981 , n1984 ); 
nor ( n1986 , n1980 , n1985 ); 
nand ( n1987 , n1940 , n1986 ); 
not ( n1988 , n1987 ); 
not ( n1989 , n1939 ); 
not ( n1990 , n1989 ); 
not ( n1991 , n1990 ); 
not ( n1992 , n1971 ); 
not ( n1993 , n1992 ); 
nor ( n1994 , n1946 , n1902 ); 
and ( n1995 , n1912 , n1994 ); 
nand ( n1996 , n1995 , n1944 ); 
nor ( n1997 , n1993 , n1996 ); 
not ( n1998 , n1997 ); 
or ( n1999 , n1991 , n1998 ); 
not ( n2000 , n1888 ); 
not ( n2001 , n2000 ); 
nand ( n2002 , n2001 , n1993 , n1929 ); 
nand ( n2003 , n1999 , n2002 ); 
nor ( n2004 , n1988 , n2003 ); 
not ( n2005 , n1930 ); 
not ( n2006 , n1940 ); 
nand ( n2007 , n2005 , n2006 ); 
nor ( n2008 , n1996 , n1955 ); 
not ( n2009 , n2008 ); 
nand ( n2010 , n1895 , n1917 ); 
nand ( n2011 , n2009 , n2010 ); 
nand ( n2012 , n2011 , n2006 ); 
not ( n2013 , n1939 ); 
not ( n2014 , n2013 ); 
nand ( n2015 , n2014 , n1950 ); 
nand ( n2016 , n2007 , n2012 , n2015 ); 
buf ( n2017 , n2000 ); 
buf ( n2018 , n2017 ); 
not ( n2019 , n2018 ); 
not ( n2020 , n1955 ); 
nand ( n2021 , n1912 , n1902 , n1966 ); 
nor ( n2022 , n1928 , n2021 ); 
nand ( n2023 , n2020 , n2022 ); 
nor ( n2024 , n2019 , n2023 ); 
nor ( n2025 , n2016 , n2024 ); 
nand ( n2026 , n1978 , n2004 , n2025 ); 
buf ( n2027 , n1943 ); 
nand ( n2028 , n2027 , n1926 ); 
not ( n2029 , n2028 ); 
nand ( n2030 , n2029 , n2020 , n2017 ); 
nor ( n2031 , n1912 , n1983 ); 
not ( n2032 , n2031 ); 
not ( n2033 , n2027 ); 
nor ( n2034 , n2032 , n2033 ); 
nand ( n2035 , n1935 , n2034 ); 
nand ( n2036 , n2030 , n2035 ); 
not ( n2037 , n2036 ); 
and ( n2038 , n1943 , n1984 ); 
nand ( n2039 , n1956 , n2038 ); 
nor ( n2040 , n2014 , n2039 ); 
not ( n2041 , n2040 ); 
not ( n2042 , n2017 ); 
nor ( n2043 , n2028 , n1942 ); 
not ( n2044 , n2043 ); 
or ( n2045 , n2042 , n2044 ); 
not ( n2046 , n1895 ); 
not ( n2047 , n1995 ); 
nor ( n2048 , n2047 , n1981 ); 
nand ( n2049 , n1989 , n2046 , n2048 ); 
nand ( n2050 , n2045 , n2049 ); 
not ( n2051 , n2050 ); 
nand ( n2052 , n2037 , n2041 , n2051 ); 
not ( n2053 , n1979 ); 
not ( n2054 , n1985 ); 
nand ( n2055 , n1890 , n2053 , n2054 ); 
not ( n2056 , n2055 ); 
not ( n2057 , n2056 ); 
not ( n2058 , n1941 ); 
nand ( n2059 , n1948 , n2058 , n1928 ); 
not ( n2060 , n2059 ); 
nand ( n2061 , n1961 , n1994 ); 
nor ( n2062 , n1981 , n2061 ); 
nand ( n2063 , n1992 , n2062 ); 
not ( n2064 , n2063 ); 
or ( n2065 , n2060 , n2064 ); 
nand ( n2066 , n2065 , n2018 ); 
nand ( n2067 , n2057 , n2066 ); 
nor ( n2068 , n2052 , n2067 ); 
not ( n2069 , n2059 ); 
nand ( n2070 , n2069 , n1922 ); 
not ( n2071 , n1895 ); 
nand ( n2072 , n2071 , n1890 , n2034 ); 
not ( n2073 , n2072 ); 
nand ( n2074 , n2043 , n2001 ); 
not ( n2075 , n2074 ); 
nor ( n2076 , n2073 , n2075 ); 
nand ( n2077 , n2070 , n2076 ); 
not ( n2078 , n2063 ); 
nand ( n2079 , n1990 , n2078 ); 
nor ( n2080 , n1928 , n2061 ); 
nand ( n2081 , n1889 , n1942 , n2080 ); 
not ( n2082 , n2081 ); 
nand ( n2083 , n2038 , n1992 ); 
nor ( n2084 , n2083 , n2013 ); 
nor ( n2085 , n2082 , n2084 ); 
nor ( n2086 , n1893 , n1915 ); 
not ( n2087 , n1913 ); 
nand ( n2088 , n2086 , n2087 ); 
not ( n2089 , n2088 ); 
nand ( n2090 , n2089 , n1922 ); 
nor ( n2091 , n2033 , n2021 ); 
nand ( n2092 , n2053 , n2091 ); 
not ( n2093 , n2092 ); 
nand ( n2094 , n2006 , n2093 ); 
nand ( n2095 , n2079 , n2085 , n2090 , n2094 ); 
nor ( n2096 , n2077 , n2095 ); 
nand ( n2097 , n2068 , n2096 ); 
nor ( n2098 , n2026 , n2097 ); 
not ( n2099 , n2098 ); 
or ( n2100 , n1882 , n2099 ); 
nand ( n2101 , n2100 , n391 ); 
not ( n2102 , n2026 ); 
and ( n2103 , n2102 , n2068 , n2096 ); 
nor ( n2104 , n2103 , n1881 ); 
or ( n2105 , n2101 , n2104 ); 
not ( n2106 , n121 ); 
or ( n2107 , n2106 , n402 ); 
nand ( n2108 , n2105 , n2107 ); 
nand ( n2109 , n1891 , n1997 ); 
nand ( n2110 , n2109 , n1951 , n2081 ); 
not ( n2111 , n1962 ); 
not ( n2112 , n2111 ); 
not ( n2113 , n2000 ); 
not ( n2114 , n1960 ); 
not ( n2115 , n1914 ); 
nand ( n2116 , n2115 , n1904 ); 
not ( n2117 , n2116 ); 
nand ( n2118 , n2113 , n2114 , n1955 , n2117 ); 
nand ( n2119 , n1888 , n1893 , n1964 ); 
not ( n2120 , n1946 ); 
nand ( n2121 , n2120 , n1914 ); 
nand ( n2122 , n2121 , n2116 ); 
not ( n2123 , n1893 ); 
not ( n2124 , n1888 ); 
nand ( n2125 , n2122 , n2123 , n2124 ); 
nand ( n2126 , n2119 , n2125 ); 
nand ( n2127 , n1960 , n2126 ); 
nand ( n2128 , n2118 , n2127 ); 
not ( n2129 , n2128 ); 
or ( n2130 , n2112 , n2129 ); 
nand ( n2131 , n2033 , n1935 , n2031 ); 
nand ( n2132 , n2130 , n2131 ); 
nor ( n2133 , n2110 , n2132 ); 
not ( n2134 , n2012 ); 
not ( n2135 , n2080 ); 
nor ( n2136 , n2013 , n1956 , n2135 ); 
not ( n2137 , n2136 ); 
nand ( n2138 , n2137 , n1987 ); 
nor ( n2139 , n2134 , n2138 ); 
nand ( n2140 , n2014 , n1919 ); 
nand ( n2141 , n2140 , n2002 ); 
not ( n2142 , n2010 ); 
nand ( n2143 , n1891 , n2142 ); 
nand ( n2144 , n1920 , n2143 ); 
nor ( n2145 , n2141 , n2144 ); 
nand ( n2146 , n2133 , n2139 , n2145 ); 
not ( n2147 , n2146 ); 
not ( n2148 , n2088 ); 
not ( n2149 , n2092 ); 
or ( n2150 , n2148 , n2149 ); 
nand ( n2151 , n2150 , n2018 ); 
nand ( n2152 , n2055 , n2151 ); 
nor ( n2153 , n1891 , n2023 ); 
not ( n2154 , n2153 ); 
nand ( n2155 , n2154 , n2066 , n2051 ); 
nor ( n2156 , n2152 , n2155 ); 
nand ( n2157 , n2001 , n2020 , n2062 ); 
not ( n2158 , n2039 ); 
nand ( n2159 , n1990 , n2158 ); 
nand ( n2160 , n2157 , n2159 , n2094 ); 
not ( n2161 , n2160 ); 
not ( n2162 , n2083 ); 
nand ( n2163 , n2018 , n2162 ); 
not ( n2164 , n2048 ); 
nor ( n2165 , n2164 , n2071 ); 
nand ( n2166 , n1990 , n2165 ); 
nand ( n2167 , n2072 , n2166 ); 
nand ( n2168 , n2070 , n2074 ); 
nor ( n2169 , n2167 , n2168 ); 
and ( n2170 , n2161 , n2163 , n2169 ); 
nand ( n2171 , n2147 , n2156 , n2170 ); 
or ( n2172 , n87 , n2171 ); 
nand ( n2173 , n2172 , n391 ); 
and ( n2174 , n2147 , n2156 , n2170 ); 
not ( n2175 , n87 ); 
nor ( n2176 , n2174 , n2175 ); 
or ( n2177 , n2173 , n2176 ); 
not ( n2178 , n96 ); 
or ( n2179 , n2178 , n402 ); 
nand ( n2180 , n2177 , n2179 ); 
and ( n2181 , n402 , n1606 ); 
not ( n2182 , n402 ); 
not ( n2183 , n134 ); 
and ( n2184 , n2182 , n2183 ); 
nor ( n2185 , n2181 , n2184 ); 
not ( n2186 , n107 ); 
not ( n2187 , n2186 ); 
nor ( n2188 , n1857 , n323 ); 
and ( n2189 , n257 , n270 ); 
nor ( n2190 , n244 , n1624 ); 
and ( n2191 , n2188 , n2189 , n2190 ); 
not ( n2192 , n325 ); 
not ( n2193 , n1670 ); 
nor ( n2194 , n2192 , n2193 ); 
not ( n2195 , n1864 ); 
nor ( n2196 , n2195 , n314 ); 
not ( n2197 , n1664 ); 
not ( n2198 , n1671 ); 
and ( n2199 , n2196 , n328 , n2197 , n2198 ); 
nand ( n2200 , n2191 , n2194 , n2199 ); 
not ( n2201 , n1852 ); 
nand ( n2202 , n2201 , n1827 , n303 ); 
not ( n2203 , n2202 ); 
not ( n2204 , n317 ); 
nand ( n2205 , n1640 , n1638 ); 
and ( n2206 , n357 , n1635 ); 
nor ( n2207 , n2206 , n284 ); 
and ( n2208 , n2205 , n2207 ); 
not ( n2209 , n1637 ); 
nand ( n2210 , n2209 , n1633 ); 
not ( n2211 , n210 ); 
nor ( n2212 , n227 , n249 ); 
and ( n2213 , n2210 , n2211 , n2212 ); 
nor ( n2214 , n2208 , n2213 ); 
or ( n2215 , n2204 , n2214 ); 
nand ( n2216 , n2215 , n1847 , n1632 ); 
nand ( n2217 , n1659 , n372 ); 
nor ( n2218 , n2216 , n2217 ); 
and ( n2219 , n363 , n1660 ); 
nand ( n2220 , n2203 , n2218 , n224 , n2219 ); 
nor ( n2221 , n2200 , n2220 ); 
not ( n2222 , n2221 ); 
or ( n2223 , n2187 , n2222 ); 
nand ( n2224 , n2223 , n402 ); 
nor ( n2225 , n2186 , n2221 ); 
or ( n2226 , n2224 , n2225 ); 
not ( n2227 , n108 ); 
or ( n2228 , n2227 , n402 ); 
nand ( n2229 , n2226 , n2228 ); 
and ( n2230 , n1 , n388 ); 
and ( n2231 , n2 , n3 ); 
nor ( n2232 , n2230 , n2231 ); 
and ( n2233 , n391 , n2232 ); 
not ( n2234 , n391 ); 
nor ( n2235 , n1495 , n1527 ); 
nand ( n2236 , n1454 , n1420 ); 
not ( n2237 , n2236 ); 
nand ( n2238 , n2235 , n1498 , n1573 , n2237 ); 
not ( n2239 , n1493 ); 
nand ( n2240 , n1497 , n1388 , n2239 ); 
not ( n2241 , n2240 ); 
nor ( n2242 , n1489 , n1456 ); 
or ( n2243 , n1395 , n2242 ); 
not ( n2244 , n1488 ); 
nand ( n2245 , n1456 , n2244 ); 
nand ( n2246 , n1395 , n2245 ); 
nand ( n2247 , n2243 , n2246 , n1540 ); 
not ( n2248 , n2247 ); 
or ( n2249 , n2241 , n2248 ); 
not ( n2250 , n1500 ); 
nor ( n2251 , n1405 , n2250 ); 
nand ( n2252 , n2249 , n2251 ); 
nand ( n2253 , n2238 , n2252 ); 
nand ( n2254 , n1450 , n1486 ); 
not ( n2255 , n1457 ); 
nand ( n2256 , n2255 , n1594 ); 
not ( n2257 , n2256 ); 
nand ( n2258 , n2257 , n1389 , n1425 ); 
not ( n2259 , n1396 ); 
nor ( n2260 , n1434 , n2259 ); 
not ( n2261 , n2260 ); 
nand ( n2262 , n2258 , n2261 ); 
nor ( n2263 , n2253 , n2254 , n2262 ); 
and ( n2264 , n1470 , n1459 ); 
nand ( n2265 , n1522 , n1589 ); 
not ( n2266 , n2265 ); 
nor ( n2267 , n2266 , n1464 ); 
nand ( n2268 , n1438 , n1586 ); 
not ( n2269 , n2268 ); 
not ( n2270 , n1423 ); 
not ( n2271 , n1517 ); 
not ( n2272 , n1451 ); 
nand ( n2273 , n2271 , n2272 , n1467 , n1558 ); 
nand ( n2274 , n2273 , n1481 ); 
nor ( n2275 , n2269 , n2270 , n2274 ); 
and ( n2276 , n2263 , n2264 , n2267 , n2275 ); 
not ( n2277 , n1542 ); 
not ( n2278 , n1472 ); 
nand ( n2279 , n2278 , n2259 , n1528 , n1501 ); 
not ( n2280 , n2279 ); 
nor ( n2281 , n2277 , n2280 ); 
not ( n2282 , n1556 ); 
nor ( n2283 , n2282 , n1569 ); 
nand ( n2284 , n1541 , n1555 ); 
nor ( n2285 , n1442 , n1509 ); 
nand ( n2286 , n1572 , n1573 , n2285 ); 
and ( n2287 , n2284 , n2286 ); 
not ( n2288 , n1547 ); 
not ( n2289 , n1565 ); 
nor ( n2290 , n2288 , n2289 ); 
nand ( n2291 , n2281 , n2283 , n2287 , n2290 ); 
and ( n2292 , n1421 , n1469 ); 
nand ( n2293 , n2292 , n1452 , n1389 ); 
nand ( n2294 , n2293 , n1580 ); 
not ( n2295 , n1555 ); 
not ( n2296 , n1582 ); 
or ( n2297 , n2295 , n2296 ); 
not ( n2298 , n1578 ); 
nand ( n2299 , n2297 , n2298 ); 
nor ( n2300 , n2294 , n2299 ); 
not ( n2301 , n1595 ); 
nor ( n2302 , n2301 , n1575 ); 
nor ( n2303 , n1452 , n1550 ); 
not ( n2304 , n2303 ); 
not ( n2305 , n2304 ); 
nand ( n2306 , n1577 , n1576 ); 
nor ( n2307 , n2306 , n1425 ); 
not ( n2308 , n2307 ); 
not ( n2309 , n2308 ); 
nor ( n2310 , n2305 , n2309 ); 
nand ( n2311 , n2300 , n2302 , n2310 ); 
nor ( n2312 , n2291 , n2311 ); 
nand ( n2313 , n2276 , n2312 ); 
not ( n2314 , n4 ); 
and ( n2315 , n2313 , n2314 ); 
not ( n2316 , n2313 ); 
and ( n2317 , n2316 , n4 ); 
nor ( n2318 , n2315 , n2317 ); 
and ( n2319 , n2234 , n2318 ); 
nor ( n2320 , n2233 , n2319 ); 
not ( n2321 , n82 ); 
and ( n2322 , n83 , n2321 ); 
not ( n2323 , n83 ); 
and ( n2324 , n2323 , n82 ); 
nor ( n2325 , n2322 , n2324 ); 
buf ( n2326 , n2325 ); 
xnor ( n2327 , n81 , n80 ); 
xor ( n2328 , n41 , n78 ); 
not ( n2329 , n2328 ); 
xor ( n2330 , n45 , n79 ); 
not ( n2331 , n2330 ); 
nand ( n2332 , n2327 , n2329 , n2331 ); 
not ( n2333 , n2332 ); 
nand ( n2334 , n2326 , n2333 ); 
not ( n2335 , n2334 ); 
xor ( n2336 , n84 , n66 ); 
not ( n2337 , n2336 ); 
and ( n2338 , n70 , n85 ); 
not ( n2339 , n70 ); 
not ( n2340 , n85 ); 
and ( n2341 , n2339 , n2340 ); 
nor ( n2342 , n2338 , n2341 ); 
buf ( n2343 , n2342 ); 
not ( n2344 , n2343 ); 
not ( n2345 , n2344 ); 
not ( n2346 , n2345 ); 
and ( n2347 , n2335 , n2337 , n2346 ); 
not ( n2348 , n2347 ); 
not ( n2349 , n2342 ); 
not ( n2350 , n2349 ); 
buf ( n2351 , n2350 ); 
not ( n2352 , n2351 ); 
not ( n2353 , n2352 ); 
buf ( n2354 , n2336 ); 
not ( n2355 , n2354 ); 
buf ( n2356 , n2325 ); 
not ( n2357 , n2356 ); 
xor ( n2358 , n80 , n81 ); 
nand ( n2359 , n2358 , n2328 , n2330 ); 
not ( n2360 , n2359 ); 
nand ( n2361 , n2357 , n2360 ); 
nor ( n2362 , n2355 , n2361 ); 
nand ( n2363 , n2353 , n2362 ); 
nand ( n2364 , n2348 , n2363 ); 
not ( n2365 , n2354 ); 
not ( n2366 , n2326 ); 
and ( n2367 , n2327 , n2328 , n2331 ); 
nand ( n2368 , n2366 , n2367 ); 
nor ( n2369 , n2365 , n2368 ); 
nand ( n2370 , n2353 , n2369 ); 
not ( n2371 , n2328 ); 
nand ( n2372 , n2371 , n2330 ); 
nor ( n2373 , n2327 , n2372 ); 
nand ( n2374 , n2326 , n2373 ); 
not ( n2375 , n2374 ); 
not ( n2376 , n2351 ); 
nand ( n2377 , n2375 , n2365 , n2376 ); 
not ( n2378 , n2344 ); 
not ( n2379 , n2329 ); 
not ( n2380 , n2379 ); 
not ( n2381 , n2336 ); 
not ( n2382 , n2331 ); 
and ( n2383 , n2382 , n2358 ); 
nand ( n2384 , n2378 , n2380 , n2381 , n2383 ); 
not ( n2385 , n2384 ); 
not ( n2386 , n2336 ); 
not ( n2387 , n2328 ); 
nor ( n2388 , n2358 , n2342 ); 
not ( n2389 , n2388 ); 
or ( n2390 , n2387 , n2389 ); 
nand ( n2391 , n2358 , n2342 ); 
or ( n2392 , n2379 , n2391 ); 
nand ( n2393 , n2390 , n2392 ); 
or ( n2394 , n2386 , n2393 ); 
buf ( n2395 , n2382 ); 
not ( n2396 , n2395 ); 
not ( n2397 , n2329 ); 
nand ( n2398 , n2397 , n2358 ); 
or ( n2399 , n2350 , n2398 ); 
not ( n2400 , n2336 ); 
nand ( n2401 , n2399 , n2400 ); 
nand ( n2402 , n2394 , n2396 , n2401 ); 
not ( n2403 , n2402 ); 
or ( n2404 , n2385 , n2403 ); 
nand ( n2405 , n2404 , n2326 ); 
nand ( n2406 , n2370 , n2377 , n2405 ); 
nor ( n2407 , n2364 , n2406 ); 
nand ( n2408 , n2386 , n2344 ); 
and ( n2409 , n2327 , n2328 , n2330 ); 
nand ( n2410 , n2326 , n2409 ); 
nor ( n2411 , n2408 , n2410 ); 
buf ( n2412 , n2345 ); 
buf ( n2413 , n2336 ); 
not ( n2414 , n2413 ); 
not ( n2415 , n2372 ); 
nand ( n2416 , n2327 , n2415 ); 
nor ( n2417 , n2326 , n2416 ); 
nand ( n2418 , n2412 , n2414 , n2417 ); 
not ( n2419 , n2351 ); 
not ( n2420 , n2356 ); 
nand ( n2421 , n2420 , n2400 , n2333 ); 
or ( n2422 , n2419 , n2421 ); 
nand ( n2423 , n2418 , n2422 ); 
nor ( n2424 , n2411 , n2423 ); 
buf ( n2425 , n2350 ); 
not ( n2426 , n2425 ); 
not ( n2427 , n2426 ); 
not ( n2428 , n2337 ); 
and ( n2429 , n2358 , n2329 , n2331 ); 
nand ( n2430 , n2357 , n2429 ); 
nor ( n2431 , n2428 , n2430 ); 
nand ( n2432 , n2427 , n2431 ); 
not ( n2433 , n2400 ); 
nand ( n2434 , n2420 , n2409 ); 
nor ( n2435 , n2433 , n2434 ); 
nand ( n2436 , n2352 , n2435 ); 
nand ( n2437 , n2381 , n2344 ); 
nor ( n2438 , n2368 , n2437 ); 
not ( n2439 , n2438 ); 
nand ( n2440 , n2436 , n2439 ); 
nor ( n2441 , n2357 , n2416 ); 
nand ( n2442 , n2351 , n2337 , n2441 ); 
not ( n2443 , n2442 ); 
not ( n2444 , n2443 ); 
nand ( n2445 , n2426 , n2431 ); 
nand ( n2446 , n2444 , n2445 ); 
nor ( n2447 , n2440 , n2446 ); 
and ( n2448 , n2407 , n2424 , n2432 , n2447 ); 
nor ( n2449 , n2355 , n2334 ); 
nand ( n2450 , n2353 , n2449 ); 
nor ( n2451 , n2420 , n2359 ); 
nand ( n2452 , n2413 , n2451 ); 
not ( n2453 , n2452 ); 
nand ( n2454 , n2353 , n2453 ); 
nor ( n2455 , n2337 , n2410 ); 
nand ( n2456 , n2412 , n2455 ); 
nand ( n2457 , n2450 , n2454 , n2456 ); 
not ( n2458 , n2457 ); 
nand ( n2459 , n2425 , n2433 , n2417 ); 
not ( n2460 , n2459 ); 
not ( n2461 , n2460 ); 
not ( n2462 , n2425 ); 
not ( n2463 , n2381 ); 
not ( n2464 , n2434 ); 
nand ( n2465 , n2462 , n2463 , n2464 ); 
nand ( n2466 , n2397 , n2331 ); 
nor ( n2467 , n2327 , n2466 ); 
not ( n2468 , n2467 ); 
nor ( n2469 , n2326 , n2468 ); 
nand ( n2470 , n2352 , n2463 , n2469 ); 
nand ( n2471 , n2461 , n2465 , n2470 ); 
not ( n2472 , n2471 ); 
buf ( n2473 , n2425 ); 
nand ( n2474 , n2366 , n2373 ); 
nor ( n2475 , n2414 , n2474 ); 
nand ( n2476 , n2473 , n2475 ); 
not ( n2477 , n2476 ); 
nor ( n2478 , n2412 , n2452 ); 
nor ( n2479 , n2477 , n2478 ); 
nand ( n2480 , n2458 , n2472 , n2479 ); 
nand ( n2481 , n2425 , n2337 , n2451 ); 
not ( n2482 , n2356 ); 
nor ( n2483 , n2482 , n2336 ); 
nand ( n2484 , n2483 , n2378 , n2467 ); 
nand ( n2485 , n2481 , n2484 ); 
not ( n2486 , n2345 ); 
nand ( n2487 , n2486 , n2428 , n2441 ); 
not ( n2488 , n2429 ); 
nor ( n2489 , n2366 , n2488 ); 
nand ( n2490 , n2376 , n2433 , n2489 ); 
nand ( n2491 , n2487 , n2490 ); 
nor ( n2492 , n2485 , n2491 ); 
not ( n2493 , n2427 ); 
nor ( n2494 , n2365 , n2374 ); 
nand ( n2495 , n2493 , n2494 ); 
nor ( n2496 , n2337 , n2430 ); 
nand ( n2497 , n2426 , n2496 ); 
buf ( n2498 , n2486 ); 
nor ( n2499 , n2433 , n2361 ); 
and ( n2500 , n2498 , n2499 ); 
not ( n2501 , n2498 ); 
nand ( n2502 , n2326 , n2367 ); 
nor ( n2503 , n2413 , n2502 ); 
and ( n2504 , n2501 , n2503 ); 
nor ( n2505 , n2500 , n2504 ); 
nand ( n2506 , n2492 , n2495 , n2497 , n2505 ); 
nor ( n2507 , n2480 , n2506 ); 
nand ( n2508 , n2448 , n2507 ); 
or ( n2509 , n77 , n2508 ); 
nand ( n2510 , n2509 , n402 ); 
and ( n2511 , n2448 , n2507 ); 
not ( n2512 , n77 ); 
nor ( n2513 , n2511 , n2512 ); 
or ( n2514 , n2510 , n2513 ); 
not ( n2515 , n86 ); 
or ( n2516 , n2515 , n402 ); 
nand ( n2517 , n2514 , n2516 ); 
not ( n2518 , n128 ); 
not ( n2519 , n2518 ); 
and ( n2520 , n542 , n723 ); 
nand ( n2521 , n2520 , n442 , n494 ); 
nand ( n2522 , n692 , n667 ); 
nor ( n2523 , n2521 , n2522 ); 
nor ( n2524 , n519 , n730 ); 
and ( n2525 , n2523 , n2524 , t_1 ); 
not ( n2526 , n2525 ); 
not ( n2527 , n658 ); 
not ( n2528 , n2527 ); 
nand ( n2529 , n447 , n749 , n553 , n575 ); 
and ( n2530 , n661 , n2529 ); 
nand ( n2531 , n2528 , n2530 , n639 , n544 ); 
not ( n2532 , n2531 ); 
nor ( n2533 , n698 , n703 ); 
not ( n2534 , n595 ); 
nor ( n2535 , n696 , n2534 ); 
nor ( n2536 , n740 , n611 ); 
and ( n2537 , n2535 , n2536 , n699 , n600 ); 
nand ( n2538 , n2532 , n589 , n2533 , n2537 ); 
nor ( n2539 , n2526 , n2538 ); 
not ( n2540 , n2539 ); 
or ( n2541 , n2519 , n2540 ); 
nand ( n2542 , n2541 , n391 ); 
nor ( n2543 , t_6 , n2518 ); 
or ( n2544 , n2542 , n2543 ); 
not ( n2545 , n129 ); 
or ( n2546 , n2545 , n391 ); 
nand ( n2547 , n2544 , n2546 ); 
nand ( n2548 , n2355 , n2489 ); 
nor ( n2549 , n2473 , n2548 ); 
and ( n2550 , n2396 , n2381 ); 
and ( n2551 , n2395 , n2354 ); 
nor ( n2552 , n2550 , n2551 ); 
or ( n2553 , n2379 , n2326 , n2358 ); 
or ( n2554 , n2357 , n2398 ); 
nand ( n2555 , n2553 , n2554 ); 
and ( n2556 , n2552 , n2376 , n2555 ); 
nor ( n2557 , n2549 , n2556 ); 
nand ( n2558 , n2557 , n2377 , n2454 , n2370 ); 
not ( n2559 , n2425 ); 
and ( n2560 , n2559 , n2503 ); 
not ( n2561 , n2559 ); 
nor ( n2562 , n2428 , n2474 ); 
and ( n2563 , n2561 , n2562 ); 
nor ( n2564 , n2560 , n2563 ); 
nor ( n2565 , n2411 , n2438 ); 
and ( n2566 , n2564 , n2565 ); 
or ( n2567 , n2498 , n2548 ); 
not ( n2568 , n2445 ); 
nor ( n2569 , n2568 , n2423 ); 
nand ( n2570 , n2566 , n2567 , n2569 ); 
nor ( n2571 , n2558 , n2570 ); 
not ( n2572 , n2502 ); 
nand ( n2573 , n2425 , n2463 , n2572 ); 
nand ( n2574 , n2476 , n2456 , n2573 ); 
not ( n2575 , n2574 ); 
not ( n2576 , n2427 ); 
nand ( n2577 , n2576 , n2455 ); 
nand ( n2578 , n2462 , n2362 ); 
nand ( n2579 , n2578 , n2470 ); 
not ( n2580 , n2486 ); 
nand ( n2581 , n2580 , n2494 ); 
nand ( n2582 , n2580 , n2496 ); 
nand ( n2583 , n2581 , n2582 ); 
nor ( n2584 , n2579 , n2583 ); 
nand ( n2585 , n2575 , n2577 , n2584 ); 
nand ( n2586 , n2580 , n2435 ); 
not ( n2587 , n2586 ); 
nor ( n2588 , n2587 , n2491 ); 
not ( n2589 , n2498 ); 
and ( n2590 , n2355 , n2469 ); 
nand ( n2591 , n2589 , n2590 ); 
nand ( n2592 , n2353 , n2503 ); 
and ( n2593 , n2481 , n2592 ); 
and ( n2594 , n2473 , n2449 ); 
not ( n2595 , n2473 ); 
and ( n2596 , n2595 , n2475 ); 
nor ( n2597 , n2594 , n2596 ); 
nand ( n2598 , n2588 , n2591 , n2593 , n2597 ); 
nor ( n2599 , n2585 , n2598 ); 
nand ( n2600 , n2571 , n2599 ); 
or ( n2601 , n126 , n2600 ); 
nand ( n2602 , n2601 , n402 ); 
and ( n2603 , n2571 , n2599 ); 
not ( n2604 , n126 ); 
nor ( n2605 , n2603 , n2604 ); 
or ( n2606 , n2602 , n2605 ); 
not ( n2607 , n127 ); 
or ( n2608 , n2607 , n402 ); 
nand ( n2609 , n2606 , n2608 ); 
not ( n2610 , n115 ); 
and ( n2611 , n1691 , n2610 ); 
not ( n2612 , n1691 ); 
and ( n2613 , n2612 , n2318 ); 
nor ( n2614 , n2611 , n2613 ); 
not ( n2615 , n2131 ); 
nor ( n2616 , n2615 , n1931 ); 
not ( n2617 , n1960 ); 
not ( n2618 , n2617 ); 
not ( n2619 , n1936 ); 
not ( n2620 , n1966 ); 
nand ( n2621 , n2619 , n2620 , n2111 ); 
not ( n2622 , n2121 ); 
not ( n2623 , n1973 ); 
not ( n2624 , n1887 ); 
nand ( n2625 , n1912 , n2624 ); 
nand ( n2626 , n2623 , n2625 ); 
nand ( n2627 , n1894 , n2622 , n2626 ); 
nand ( n2628 , n2621 , n2627 ); 
not ( n2629 , n2628 ); 
or ( n2630 , n2618 , n2629 ); 
nand ( n2631 , n2630 , n1958 ); 
not ( n2632 , n1983 ); 
nand ( n2633 , n1928 , n1992 , n2632 , n1973 ); 
nand ( n2634 , n2633 , n2081 ); 
nor ( n2635 , n2631 , n2634 ); 
and ( n2636 , n2616 , n2635 ); 
nand ( n2637 , n2140 , n2015 ); 
nor ( n2638 , n2637 , n2003 ); 
nand ( n2639 , n1935 , n2022 ); 
nand ( n2640 , n2639 , n2143 ); 
nor ( n2641 , n2138 , n2640 ); 
and ( n2642 , n2636 , n2638 , n2641 ); 
nand ( n2643 , n2018 , n2165 ); 
not ( n2644 , n2001 ); 
not ( n2645 , n1986 ); 
or ( n2646 , n2644 , n2645 ); 
nand ( n2647 , n2646 , n2055 ); 
not ( n2648 , n2647 ); 
nand ( n2649 , n2643 , n2066 , n2648 ); 
nand ( n2650 , n2030 , n2151 ); 
nor ( n2651 , n2649 , n2650 ); 
not ( n2652 , n2084 ); 
nand ( n2653 , n2001 , n1993 , n2091 ); 
nand ( n2654 , n2652 , n2090 , n2653 ); 
not ( n2655 , n2654 ); 
not ( n2656 , n2157 ); 
nor ( n2657 , n2656 , n2040 ); 
and ( n2658 , n2655 , n2657 , n2166 , n2076 ); 
and ( n2659 , n2642 , n2651 , n2658 ); 
not ( n2660 , n130 ); 
nor ( n2661 , n2659 , n2660 ); 
nand ( n2662 , n2642 , n2651 , n2658 ); 
or ( n2663 , n2662 , n130 ); 
nand ( n2664 , n2663 , n391 ); 
or ( n2665 , n2661 , n2664 ); 
not ( n2666 , n131 ); 
or ( n2667 , n2666 , n402 ); 
nand ( n2668 , n2665 , n2667 ); 
not ( n2669 , n2280 ); 
nor ( n2670 , n1454 , n1420 ); 
not ( n2671 , n2670 ); 
nand ( n2672 , n2671 , n2236 ); 
and ( n2673 , n1506 , n2672 ); 
nor ( n2674 , n1507 , n1404 , n1479 ); 
nor ( n2675 , n2673 , n2674 ); 
or ( n2676 , n1495 , n2675 ); 
not ( n2677 , n1533 ); 
nor ( n2678 , n1420 , n1479 ); 
nand ( n2679 , n2677 , n2678 ); 
nand ( n2680 , n2676 , n2679 ); 
and ( n2681 , n2680 , n1505 , n1499 ); 
not ( n2682 , n1448 ); 
and ( n2683 , n1576 , n2682 , n1451 ); 
nor ( n2684 , n2681 , n2683 ); 
nand ( n2685 , n2669 , n2684 , n1530 , n2286 ); 
and ( n2686 , n2258 , n1486 ); 
not ( n2687 , n1463 ); 
nor ( n2688 , n2687 , n1520 ); 
not ( n2689 , n1470 ); 
not ( n2690 , n2273 ); 
nor ( n2691 , n2689 , n2690 ); 
and ( n2692 , n2691 , n1441 , n2268 ); 
nand ( n2693 , n2686 , n2688 , n2692 ); 
nor ( n2694 , n2685 , n2693 ); 
and ( n2695 , n1568 , n1545 ); 
and ( n2696 , n1522 , n1567 ); 
nor ( n2697 , n1557 , n2696 ); 
not ( n2698 , n1562 ); 
nor ( n2699 , n1389 , n2256 ); 
nand ( n2700 , n1515 , n2699 ); 
not ( n2701 , n2700 ); 
nor ( n2702 , n2701 , n1553 ); 
and ( n2703 , n2695 , n2697 , n2698 , n2702 ); 
not ( n2704 , n2294 ); 
and ( n2705 , n1388 , n1451 , n1421 , n1510 ); 
not ( n2706 , n2705 ); 
nand ( n2707 , n2706 , n1590 ); 
not ( n2708 , n2303 ); 
nand ( n2709 , n2708 , n2308 ); 
nor ( n2710 , n2707 , n2709 ); 
nand ( n2711 , n2704 , n2710 , n1598 ); 
not ( n2712 , n2711 ); 
nand ( n2713 , n2694 , n2703 , n2712 ); 
or ( n2714 , n2713 , n75 ); 
nand ( n2715 , n2714 , n391 ); 
and ( n2716 , n2694 , n2703 , n2712 ); 
not ( n2717 , n75 ); 
nor ( n2718 , n2716 , n2717 ); 
or ( n2719 , n2715 , n2718 ); 
not ( n2720 , n76 ); 
or ( n2721 , n2720 , n402 ); 
nand ( n2722 , n2719 , n2721 ); 
nor ( n2723 , n2549 , n2347 ); 
not ( n2724 , n2326 ); 
not ( n2725 , n2395 ); 
nand ( n2726 , n2358 , n2379 , n2343 ); 
not ( n2727 , n2726 ); 
and ( n2728 , n2725 , n2727 ); 
not ( n2729 , n2397 ); 
nand ( n2730 , n2729 , n2349 ); 
nor ( n2731 , n2358 , n2730 ); 
and ( n2732 , n2395 , n2731 ); 
nor ( n2733 , n2728 , n2732 ); 
or ( n2734 , n2414 , n2733 ); 
nand ( n2735 , n2397 , n2343 ); 
not ( n2736 , n2735 ); 
not ( n2737 , n2730 ); 
or ( n2738 , n2736 , n2737 ); 
nand ( n2739 , n2738 , n2383 ); 
or ( n2740 , n2463 , n2739 ); 
nand ( n2741 , n2734 , n2740 ); 
nand ( n2742 , n2724 , n2741 ); 
nand ( n2743 , n2723 , n2742 , n2363 , n2456 ); 
and ( n2744 , n2377 , n2564 ); 
not ( n2745 , n2427 ); 
not ( n2746 , n2421 ); 
nand ( n2747 , n2745 , n2746 ); 
nand ( n2748 , n2442 , n2422 ); 
not ( n2749 , n2436 ); 
nor ( n2750 , n2748 , n2749 , n2411 ); 
nand ( n2751 , n2744 , n2747 , n2750 ); 
nor ( n2752 , n2743 , n2751 ); 
nand ( n2753 , n2470 , n2581 , n2459 ); 
not ( n2754 , n2753 ); 
not ( n2755 , n2427 ); 
nand ( n2756 , n2755 , n2369 ); 
not ( n2757 , n2478 ); 
nand ( n2758 , n2757 , n2582 ); 
nand ( n2759 , n2578 , n2573 ); 
nor ( n2760 , n2758 , n2759 ); 
nand ( n2761 , n2754 , n2756 , n2760 ); 
not ( n2762 , n2484 ); 
not ( n2763 , n2462 ); 
not ( n2764 , n2449 ); 
or ( n2765 , n2763 , n2764 ); 
nand ( n2766 , n2765 , n2487 ); 
nor ( n2767 , n2762 , n2766 ); 
nand ( n2768 , n2498 , n2590 ); 
and ( n2769 , n2481 , n2586 ); 
and ( n2770 , n2497 , n2490 ); 
nand ( n2771 , n2767 , n2768 , n2769 , n2770 ); 
nor ( n2772 , n2761 , n2771 ); 
nand ( n2773 , n2752 , n2772 ); 
or ( n2774 , n116 , n2773 ); 
nand ( n2775 , n2774 , n391 ); 
and ( n2776 , n2752 , n2772 ); 
not ( n2777 , n116 ); 
nor ( n2778 , n2776 , n2777 ); 
or ( n2779 , n2775 , n2778 ); 
not ( n2780 , n117 ); 
or ( n2781 , n2780 , n402 ); 
nand ( n2782 , n2779 , n2781 ); 
not ( n2783 , n830 ); 
and ( n2784 , n877 , n818 ); 
not ( n2785 , n809 ); 
not ( n2786 , n826 ); 
or ( n2787 , n2785 , n2786 ); 
nand ( n2788 , n2787 , n1703 ); 
nand ( n2789 , n845 , n2788 ); 
nor ( n2790 , n2784 , n2789 ); 
nor ( n2791 , n2783 , n2790 ); 
and ( n2792 , n2791 , n932 , n937 , n949 ); 
not ( n2793 , n979 ); 
nand ( n2794 , n2793 , n854 ); 
not ( n2795 , n1033 ); 
nand ( n2796 , n2795 , n1036 ); 
nor ( n2797 , n2794 , n2796 ); 
and ( n2798 , n2792 , n2797 , n994 , n1716 ); 
nor ( n2799 , n921 , n1063 ); 
not ( n2800 , n1726 ); 
and ( n2801 , n2799 , n1725 , n1060 , n2800 ); 
nor ( n2802 , n875 , n1053 ); 
not ( n2803 , n1733 ); 
not ( n2804 , n1737 ); 
nor ( n2805 , n2804 , n1056 ); 
and ( n2806 , n2802 , n2803 , n2805 ); 
nand ( n2807 , n2798 , n2801 , n2806 ); 
or ( n2808 , n124 , n2807 ); 
nand ( n2809 , n2808 , n402 ); 
and ( n2810 , n2798 , n2801 , n2806 ); 
not ( n2811 , n124 ); 
nor ( n2812 , n2810 , n2811 ); 
or ( n2813 , n2809 , n2812 ); 
not ( n2814 , n125 ); 
or ( n2815 , n2814 , n402 ); 
nand ( n2816 , n2813 , n2815 ); 
nor ( n2817 , n2705 , n1435 ); 
not ( n2818 , n2274 ); 
nand ( n2819 , n2817 , n2265 , n2818 ); 
not ( n2820 , n2819 ); 
nor ( n2821 , n1499 , n1396 , n2679 ); 
nor ( n2822 , n2821 , n1487 ); 
nor ( n2823 , n2260 , n2683 ); 
not ( n2824 , n1502 ); 
nor ( n2825 , n1497 , n1428 ); 
not ( n2826 , n1466 ); 
nand ( n2827 , n2825 , n2826 , n2239 ); 
not ( n2828 , n1394 ); 
nor ( n2829 , n1387 , n2828 ); 
not ( n2830 , n1405 ); 
not ( n2831 , n1454 ); 
or ( n2832 , n2830 , n2831 ); 
or ( n2833 , n1454 , n1405 ); 
nand ( n2834 , n2832 , n2833 ); 
nand ( n2835 , n2829 , n1497 , n2834 ); 
nand ( n2836 , n2827 , n2835 ); 
nand ( n2837 , n2824 , n2836 ); 
and ( n2838 , n1530 , n2822 , n2823 , n2837 ); 
not ( n2839 , n1459 ); 
nor ( n2840 , n2839 , n1591 ); 
nand ( n2841 , n2820 , n2838 , n2840 ); 
and ( n2842 , n1514 , n1511 ); 
not ( n2843 , n1514 ); 
and ( n2844 , n2843 , n1567 ); 
nor ( n2845 , n2842 , n2844 ); 
nand ( n2846 , n2845 , n2284 , n1565 ); 
nand ( n2847 , n2279 , n1552 ); 
nor ( n2848 , n2846 , n2847 ); 
nor ( n2849 , n2294 , n2299 ); 
nand ( n2850 , n1583 , n2700 ); 
not ( n2851 , n2307 ); 
nand ( n2852 , n2851 , n1595 ); 
nor ( n2853 , n2850 , n2852 ); 
nand ( n2854 , n2848 , n2849 , n2853 , n2695 ); 
nor ( n2855 , n2841 , n2854 ); 
not ( n2856 , n2855 ); 
not ( n2857 , n55 ); 
and ( n2858 , n2856 , n2857 ); 
nor ( n2859 , n2841 , n2854 ); 
and ( n2860 , n55 , n2859 ); 
nor ( n2861 , n2858 , n2860 ); 
and ( n2862 , n391 , n2861 ); 
not ( n2863 , n391 ); 
not ( n2864 , n109 ); 
and ( n2865 , n2863 , n2864 ); 
nor ( n2866 , n2862 , n2865 ); 
and ( n2867 , n54 , n388 ); 
and ( n2868 , n3 , n35 ); 
nor ( n2869 , n2867 , n2868 ); 
and ( n2870 , n391 , n2869 ); 
not ( n2871 , n391 ); 
and ( n2872 , n2871 , n2861 ); 
nor ( n2873 , n2870 , n2872 ); 
patch p0 (.t_0(t_0), .t_1(t_1), .t_2(t_2), .t_3(t_3), .t_4(t_4), .t_5(t_5), .t_6(t_6), .t_7(t_7), .g1(n708), .g2(n420), .g3(n414), .g4(n423), .g5(n437), .g6(n644), .g7(n434), .g8(n454), .g9(n456), .g10(n407), .g11(n390), .g12(n719), .g13(n2519));
endmodule 

