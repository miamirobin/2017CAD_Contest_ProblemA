module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 ; 
output g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 ; 
wire t_0 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( n158 , g157 ); 
buf ( n159 , g158 ); 
buf ( n160 , g159 ); 
buf ( n161 , g160 ); 
buf ( n162 , g161 ); 
buf ( n163 , g162 ); 
buf ( n164 , g163 ); 
buf ( n165 , g164 ); 
buf ( n166 , g165 ); 
buf ( n167 , g166 ); 
buf ( n168 , g167 ); 
buf ( n169 , g168 ); 
buf ( n170 , g169 ); 
buf ( n171 , g170 ); 
buf ( n172 , g171 ); 
buf ( n173 , g172 ); 
buf ( n174 , g173 ); 
buf ( n175 , g174 ); 
buf ( n176 , g175 ); 
buf ( n177 , g176 ); 
buf ( n178 , g177 ); 
buf ( n179 , g178 ); 
buf ( n180 , g179 ); 
buf ( n181 , g180 ); 
buf ( n182 , g181 ); 
buf ( n183 , g182 ); 
buf ( n184 , g183 ); 
buf ( n185 , g184 ); 
buf ( n186 , g185 ); 
buf ( n187 , g186 ); 
buf ( n188 , g187 ); 
buf ( n189 , g188 ); 
buf ( n190 , g189 ); 
buf ( n191 , g190 ); 
buf ( n192 , g191 ); 
buf ( n193 , g192 ); 
buf ( n194 , g193 ); 
buf ( n195 , g194 ); 
buf ( n196 , g195 ); 
buf ( n197 , g196 ); 
buf ( n198 , g197 ); 
buf ( n199 , g198 ); 
buf ( n200 , g199 ); 
buf ( n201 , g200 ); 
buf ( n202 , g201 ); 
buf ( n203 , g202 ); 
buf ( n204 , g203 ); 
buf ( n205 , g204 ); 
buf ( n206 , g205 ); 
buf ( n207 , g206 ); 
buf ( n208 , g207 ); 
buf ( n209 , g208 ); 
buf ( n210 , g209 ); 
buf ( n211 , g210 ); 
buf ( n212 , g211 ); 
buf ( n213 , g212 ); 
buf ( n214 , g213 ); 
buf ( n215 , g214 ); 
buf ( n216 , g215 ); 
buf ( n217 , g216 ); 
buf ( n218 , g217 ); 
buf ( n219 , g218 ); 
buf ( n220 , g219 ); 
buf ( n221 , g220 ); 
buf ( n222 , g221 ); 
buf ( n223 , g222 ); 
buf ( n224 , g223 ); 
buf ( n225 , g224 ); 
buf ( n226 , g225 ); 
buf ( n227 , g226 ); 
buf ( n228 , g227 ); 
buf ( n229 , g228 ); 
buf ( n230 , g229 ); 
buf ( n231 , g230 ); 
buf ( n232 , g231 ); 
buf ( n233 , g232 ); 
buf ( n234 , g233 ); 
buf ( n235 , g234 ); 
buf ( n236 , g235 ); 
buf ( n237 , g236 ); 
buf ( n238 , g237 ); 
buf ( n239 , g238 ); 
buf ( n240 , g239 ); 
buf ( n241 , g240 ); 
buf ( n242 , g241 ); 
buf ( n243 , g242 ); 
buf ( n244 , g243 ); 
buf ( n245 , g244 ); 
buf ( n246 , g245 ); 
buf ( n247 , g246 ); 
buf ( n248 , g247 ); 
buf ( n249 , g248 ); 
buf ( n250 , g249 ); 
buf ( n251 , g250 ); 
buf ( n252 , g251 ); 
buf ( n253 , g252 ); 
buf ( n254 , g253 ); 
buf ( n255 , g254 ); 
buf ( n256 , g255 ); 
buf ( n257 , g256 ); 
buf ( n258 , g257 ); 
buf ( n259 , g258 ); 
buf ( n260 , g259 ); 
buf ( n261 , g260 ); 
buf ( n262 , g261 ); 
buf ( n263 , g262 ); 
buf ( n264 , g263 ); 
buf ( n265 , g264 ); 
buf ( n266 , g265 ); 
buf ( n267 , g266 ); 
buf ( n268 , g267 ); 
buf ( n269 , g268 ); 
buf ( n270 , g269 ); 
buf ( n271 , g270 ); 
buf ( n272 , g271 ); 
buf ( n273 , g272 ); 
buf ( n274 , g273 ); 
buf ( n275 , g274 ); 
buf ( n276 , g275 ); 
buf ( n277 , g276 ); 
buf ( n278 , g277 ); 
buf ( n279 , g278 ); 
buf ( n280 , g279 ); 
buf ( n281 , g280 ); 
buf ( n282 , g281 ); 
buf ( n283 , g282 ); 
buf ( n284 , g283 ); 
buf ( n285 , g284 ); 
buf ( n286 , g285 ); 
buf ( n287 , g286 ); 
buf ( n288 , g287 ); 
buf ( n289 , g288 ); 
buf ( n290 , g289 ); 
buf ( n291 , g290 ); 
buf ( n292 , g291 ); 
buf ( n293 , g292 ); 
buf ( n294 , g293 ); 
buf ( n295 , g294 ); 
buf ( n296 , g295 ); 
buf ( n297 , g296 ); 
buf ( n298 , g297 ); 
buf ( n299 , g298 ); 
buf ( n300 , g299 ); 
buf ( n301 , g300 ); 
buf ( n302 , g301 ); 
buf ( n303 , g302 ); 
buf ( n304 , g303 ); 
buf ( n305 , g304 ); 
buf ( n306 , g305 ); 
buf ( n307 , g306 ); 
buf ( n308 , g307 ); 
buf ( n309 , g308 ); 
buf ( n310 , g309 ); 
buf ( n311 , g310 ); 
buf ( n312 , g311 ); 
buf ( n313 , g312 ); 
buf ( n314 , g313 ); 
buf ( n315 , g314 ); 
buf ( n316 , g315 ); 
buf ( n317 , g316 ); 
buf ( n318 , g317 ); 
buf ( n319 , g318 ); 
buf ( n320 , g319 ); 
buf ( n321 , g320 ); 
buf ( n322 , g321 ); 
buf ( n323 , g322 ); 
buf ( n324 , g323 ); 
buf ( n325 , g324 ); 
buf ( n326 , g325 ); 
buf ( n327 , g326 ); 
buf ( n328 , g327 ); 
buf ( n329 , g328 ); 
buf ( n330 , g329 ); 
buf ( n331 , g330 ); 
buf ( n332 , g331 ); 
buf ( n333 , g332 ); 
buf ( n334 , g333 ); 
buf ( n335 , g334 ); 
buf ( n336 , g335 ); 
buf ( n337 , g336 ); 
buf ( n338 , g337 ); 
buf ( n339 , g338 ); 
buf ( n340 , g339 ); 
buf ( n341 , g340 ); 
buf ( n342 , g341 ); 
buf ( n343 , g342 ); 
buf ( n344 , g343 ); 
buf ( n345 , g344 ); 
buf ( n346 , g345 ); 
buf ( n347 , g346 ); 
buf ( n348 , g347 ); 
buf ( n349 , g348 ); 
buf ( n350 , g349 ); 
buf ( n351 , g350 ); 
buf ( n352 , g351 ); 
buf ( n353 , g352 ); 
buf ( n354 , g353 ); 
buf ( n355 , g354 ); 
buf ( n356 , g355 ); 
buf ( n357 , g356 ); 
buf ( n358 , g357 ); 
buf ( n359 , g358 ); 
buf ( n360 , g359 ); 
buf ( n361 , g360 ); 
buf ( n362 , g361 ); 
buf ( n363 , g362 ); 
buf ( n364 , g363 ); 
buf ( n365 , g364 ); 
buf ( n366 , g365 ); 
buf ( n367 , g366 ); 
buf ( n368 , g367 ); 
buf ( n369 , g368 ); 
buf ( n370 , g369 ); 
buf ( n371 , g370 ); 
buf ( n372 , g371 ); 
buf ( n373 , g372 ); 
buf ( n374 , g373 ); 
buf ( n375 , g374 ); 
buf ( n376 , g375 ); 
buf ( n377 , g376 ); 
buf ( n378 , g377 ); 
buf ( n379 , g378 ); 
buf ( n380 , g379 ); 
buf ( n381 , g380 ); 
buf ( n382 , g381 ); 
buf ( n383 , g382 ); 
buf ( n384 , g383 ); 
buf ( n385 , g384 ); 
buf ( n386 , g385 ); 
buf ( n387 , g386 ); 
buf ( n388 , g387 ); 
buf ( n389 , g388 ); 
buf ( n390 , g389 ); 
buf ( n391 , g390 ); 
buf ( n392 , g391 ); 
buf ( n393 , g392 ); 
buf ( n394 , g393 ); 
buf ( n395 , g394 ); 
buf ( n396 , g395 ); 
buf ( n397 , g396 ); 
buf ( n398 , g397 ); 
buf ( n399 , g398 ); 
buf ( n400 , g399 ); 
buf ( n401 , g400 ); 
buf ( n402 , g401 ); 
buf ( n403 , g402 ); 
buf ( n404 , g403 ); 
buf ( n405 , g404 ); 
buf ( n406 , g405 ); 
buf ( n407 , g406 ); 
buf ( n408 , g407 ); 
buf ( n409 , g408 ); 
buf ( n410 , g409 ); 
buf ( n411 , g410 ); 
buf ( g411 , n412 ); 
buf ( g412 , n413 ); 
buf ( g413 , n414 ); 
buf ( g414 , n415 ); 
buf ( g415 , n416 ); 
buf ( g416 , n417 ); 
buf ( g417 , n418 ); 
buf ( g418 , n419 ); 
buf ( g419 , n420 ); 
buf ( g420 , n421 ); 
buf ( g421 , n422 ); 
buf ( g422 , n423 ); 
buf ( g423 , n424 ); 
buf ( g424 , n425 ); 
buf ( g425 , n426 ); 
buf ( g426 , n427 ); 
buf ( g427 , n428 ); 
buf ( g428 , n429 ); 
buf ( g429 , n430 ); 
buf ( g430 , n431 ); 
buf ( g431 , n432 ); 
buf ( g432 , n433 ); 
buf ( g433 , n434 ); 
buf ( g434 , n435 ); 
buf ( g435 , n436 ); 
buf ( g436 , n437 ); 
buf ( g437 , n438 ); 
buf ( g438 , n439 ); 
buf ( g439 , n440 ); 
buf ( g440 , n441 ); 
buf ( g441 , n442 ); 
buf ( g442 , n443 ); 
buf ( g443 , n444 ); 
buf ( g444 , n445 ); 
buf ( g445 , n446 ); 
buf ( g446 , n447 ); 
buf ( g447 , n448 ); 
buf ( g448 , n449 ); 
buf ( g449 , n450 ); 
buf ( g450 , n451 ); 
buf ( g451 , n452 ); 
buf ( g452 , n453 ); 
buf ( g453 , n454 ); 
buf ( g454 , n455 ); 
buf ( g455 , n456 ); 
buf ( g456 , n457 ); 
buf ( g457 , n458 ); 
buf ( g458 , n459 ); 
buf ( g459 , n460 ); 
buf ( g460 , n461 ); 
buf ( g461 , n462 ); 
buf ( g462 , n463 ); 
buf ( g463 , n464 ); 
buf ( g464 , n465 ); 
buf ( g465 , n466 ); 
buf ( g466 , n467 ); 
buf ( g467 , n468 ); 
buf ( g468 , n469 ); 
buf ( g469 , n470 ); 
buf ( g470 , n471 ); 
buf ( g471 , n472 ); 
buf ( g472 , n473 ); 
buf ( g473 , n474 ); 
buf ( g474 , n475 ); 
buf ( g475 , n476 ); 
buf ( g476 , n477 ); 
buf ( g477 , n478 ); 
buf ( g478 , n479 ); 
buf ( g479 , n480 ); 
buf ( g480 , n481 ); 
buf ( g481 , n482 ); 
buf ( g482 , n483 ); 
buf ( g483 , n484 ); 
buf ( g484 , n485 ); 
buf ( g485 , n486 ); 
buf ( g486 , n487 ); 
buf ( g487 , n488 ); 
buf ( g488 , n489 ); 
buf ( g489 , n490 ); 
buf ( g490 , n491 ); 
buf ( g491 , n492 ); 
buf ( g492 , n493 ); 
buf ( g493 , n494 ); 
buf ( g494 , n495 ); 
buf ( g495 , n496 ); 
buf ( g496 , n497 ); 
buf ( g497 , n498 ); 
buf ( g498 , n499 ); 
buf ( g499 , n500 ); 
buf ( g500 , n501 ); 
buf ( g501 , n502 ); 
buf ( g502 , n503 ); 
buf ( g503 , n504 ); 
buf ( g504 , n505 ); 
buf ( g505 , n506 ); 
buf ( g506 , n507 ); 
buf ( g507 , n508 ); 
buf ( g508 , n509 ); 
buf ( g509 , n510 ); 
buf ( g510 , n511 ); 
buf ( g511 , n512 ); 
buf ( g512 , n513 ); 
buf ( g513 , n514 ); 
buf ( g514 , n515 ); 
buf ( g515 , n516 ); 
buf ( g516 , n517 ); 
buf ( g517 , n518 ); 
buf ( g518 , n519 ); 
buf ( g519 , n520 ); 
buf ( g520 , n521 ); 
buf ( g521 , n522 ); 
buf ( g522 , n523 ); 
buf ( g523 , n524 ); 
buf ( g524 , n525 ); 
buf ( g525 , n526 ); 
buf ( g526 , n527 ); 
buf ( g527 , n528 ); 
buf ( g528 , n529 ); 
buf ( g529 , n530 ); 
buf ( g530 , n531 ); 
buf ( g531 , n532 ); 
buf ( g532 , n533 ); 
buf ( g533 , n534 ); 
buf ( g534 , n535 ); 
buf ( g535 , n536 ); 
buf ( g536 , n537 ); 
buf ( g537 , n538 ); 
buf ( g538 , n539 ); 
buf ( n412 , n1030 ); 
buf ( n413 , n1603 ); 
buf ( n414 , n884 ); 
buf ( n415 , n917 ); 
buf ( n416 , n951 ); 
buf ( n417 , n983 ); 
buf ( n418 , n850 ); 
buf ( n419 , n1078 ); 
buf ( n420 , n1120 ); 
buf ( n421 , n1151 ); 
buf ( n422 , n1185 ); 
buf ( n423 , n1851 ); 
buf ( n424 , n1855 ); 
buf ( n425 , n1231 ); 
buf ( n426 , n1478 ); 
buf ( n427 , n1299 ); 
buf ( n428 , n1635 ); 
buf ( n429 , n1733 ); 
buf ( n430 , n1701 ); 
buf ( n431 , n1667 ); 
buf ( n432 , n1268 ); 
buf ( n433 , n1558 ); 
buf ( n434 , n1511 ); 
buf ( n435 , n1333 ); 
buf ( n436 , n1765 ); 
buf ( n437 , n1367 ); 
buf ( n438 , n1403 ); 
buf ( n439 , n1445 ); 
buf ( n440 , n1847 ); 
buf ( n441 , n1843 ); 
buf ( n442 , n1860 ); 
buf ( n443 , n1810 ); 
buf ( n444 , n1815 ); 
buf ( n445 , n1864 ); 
buf ( n446 , n1799 ); 
buf ( n447 , n1517 ); 
buf ( n448 , n1825 ); 
buf ( n449 , n1833 ); 
buf ( n450 , n748 ); 
buf ( n451 , n1781 ); 
buf ( n452 , n1527 ); 
buf ( n453 , n1775 ); 
buf ( n454 , n1805 ); 
buf ( n455 , n1563 ); 
buf ( n456 , n707 ); 
buf ( n457 , n1867 ); 
buf ( n458 , n1944 ); 
buf ( n459 , n16 ); 
buf ( n460 , n16 ); 
buf ( n461 , n16 ); 
buf ( n462 , n16 ); 
buf ( n463 , n16 ); 
buf ( n464 , n16 ); 
buf ( n465 , n16 ); 
buf ( n466 , n16 ); 
buf ( n467 , n16 ); 
buf ( n468 , n16 ); 
buf ( n469 , n16 ); 
buf ( n470 , n16 ); 
buf ( n471 , n16 ); 
buf ( n472 , n16 ); 
buf ( n473 , n16 ); 
buf ( n474 , n16 ); 
buf ( n475 , n16 ); 
buf ( n476 , n16 ); 
buf ( n477 , n16 ); 
buf ( n478 , n16 ); 
buf ( n479 , n16 ); 
buf ( n480 , n16 ); 
buf ( n481 , n16 ); 
buf ( n482 , n16 ); 
buf ( n483 , n16 ); 
buf ( n484 , n16 ); 
buf ( n485 , n16 ); 
buf ( n486 , n16 ); 
buf ( n487 , n16 ); 
buf ( n488 , n16 ); 
buf ( n489 , n1873 ); 
buf ( n490 , n16 ); 
buf ( n491 , n16 ); 
buf ( n492 , n1871 ); 
buf ( n493 , n16 ); 
buf ( n494 , n16 ); 
buf ( n495 , n16 ); 
buf ( n496 , n16 ); 
buf ( n497 , n16 ); 
buf ( n498 , n16 ); 
buf ( n499 , n16 ); 
buf ( n500 , n16 ); 
buf ( n501 , n1044 ); 
buf ( n502 , n1044 ); 
buf ( n503 , n1946 ); 
buf ( n504 , n16 ); 
buf ( n505 , n1947 ); 
buf ( n506 , n16 ); 
buf ( n507 , n1942 ); 
buf ( n508 , n16 ); 
buf ( n509 , n1945 ); 
buf ( n510 , n16 ); 
buf ( n511 , n16 ); 
buf ( n512 , n16 ); 
buf ( n513 , n16 ); 
buf ( n514 , n1948 ); 
buf ( n515 , n16 ); 
buf ( n516 , n16 ); 
buf ( n517 , n16 ); 
buf ( n518 , n16 ); 
buf ( n519 , n16 ); 
buf ( n520 , n544 ); 
buf ( n521 , n16 ); 
buf ( n522 , n16 ); 
buf ( n523 , n1881 ); 
buf ( n524 , n1901 ); 
buf ( n525 , n1877 ); 
buf ( n526 , n1893 ); 
buf ( n527 , n1921 ); 
buf ( n528 , n1885 ); 
buf ( n529 , n1897 ); 
buf ( n530 , n1925 ); 
buf ( n531 , n1909 ); 
buf ( n532 , n1889 ); 
buf ( n533 , n1941 ); 
buf ( n534 , n1917 ); 
buf ( n535 , n1913 ); 
buf ( n536 , n1905 ); 
buf ( n537 , n1929 ); 
buf ( n538 , n1937 ); 
buf ( n539 , n1933 ); 
and ( n544 , n371 , n348 , n370 ); 
not ( n545 , n544 ); 
nand ( n546 , n545 , n372 , n370 ); 
not ( n547 , n161 ); 
not ( n548 , n47 ); 
not ( n549 , n351 ); 
nor ( n550 , n16 , n290 ); 
nor ( n551 , n549 , n550 ); 
not ( n552 , n551 ); 
nand ( n553 , n548 , n552 ); 
not ( n554 , n550 ); 
not ( n555 , n554 ); 
nand ( n556 , n555 , n552 ); 
not ( n557 , n550 ); 
nand ( n558 , n557 , n47 , n551 ); 
nand ( n559 , n553 , n556 , n558 ); 
not ( n560 , n95 ); 
not ( n561 , n350 ); 
nor ( n562 , n16 , n245 ); 
nor ( n563 , n561 , n562 ); 
not ( n564 , n563 ); 
nand ( n565 , n560 , n564 ); 
not ( n566 , n562 ); 
not ( n567 , n566 ); 
nand ( n568 , n567 , n564 ); 
not ( n569 , n562 ); 
nand ( n570 , n569 , n95 , n563 ); 
nand ( n571 , n565 , n568 , n570 ); 
not ( n572 , n352 ); 
nor ( n573 , n16 , n318 ); 
nor ( n574 , n572 , n573 ); 
or ( n575 , n83 , n574 ); 
not ( n576 , n573 ); 
not ( n577 , n576 ); 
not ( n578 , n574 ); 
nand ( n579 , n577 , n578 ); 
not ( n580 , n573 ); 
nand ( n581 , n580 , n83 , n574 ); 
nand ( n582 , n575 , n579 , n581 ); 
nand ( n583 , n559 , n571 , n582 ); 
not ( n584 , n583 ); 
not ( n585 , n71 ); 
nor ( n586 , n16 , n195 ); 
not ( n587 , n586 ); 
nand ( n588 , n587 , n359 ); 
nand ( n589 , n585 , n588 ); 
not ( n590 , n586 ); 
not ( n591 , n590 ); 
nand ( n592 , n591 , n588 ); 
not ( n593 , n588 ); 
not ( n594 , n590 ); 
not ( n595 , n594 ); 
nand ( n596 , n593 , n595 , n71 ); 
nand ( n597 , n589 , n592 , n596 ); 
not ( n598 , n59 ); 
nor ( n599 , n16 , n306 ); 
not ( n600 , n599 ); 
nand ( n601 , n600 , n353 ); 
nand ( n602 , n598 , n601 ); 
not ( n603 , n599 ); 
not ( n604 , n603 ); 
nand ( n605 , n604 , n601 ); 
not ( n606 , n603 ); 
not ( n607 , n606 ); 
not ( n608 , n601 ); 
nand ( n609 , n607 , n59 , n608 ); 
nand ( n610 , n602 , n605 , n609 ); 
nand ( n611 , n597 , n610 ); 
not ( n612 , n611 ); 
not ( n613 , n10 ); 
not ( n614 , n356 ); 
nor ( n615 , n16 , n233 ); 
or ( n616 , n614 , n615 ); 
nand ( n617 , n613 , n616 ); 
not ( n618 , n615 ); 
not ( n619 , n618 ); 
nand ( n620 , n619 , n616 ); 
not ( n621 , n618 ); 
not ( n622 , n621 ); 
and ( n623 , n356 , n618 ); 
nand ( n624 , n622 , n10 , n623 ); 
nand ( n625 , n617 , n620 , n624 ); 
not ( n626 , n368 ); 
nor ( n627 , n16 , n283 ); 
not ( n628 , n627 ); 
nand ( n629 , n354 , n628 ); 
nand ( n630 , n626 , n629 ); 
not ( n631 , n628 ); 
nand ( n632 , n631 , n629 ); 
not ( n633 , n627 ); 
not ( n634 , n354 ); 
nor ( n635 , n634 , n627 ); 
nand ( n636 , n633 , n368 , n635 ); 
nand ( n637 , n630 , n632 , n636 ); 
and ( n638 , n625 , n637 ); 
not ( n639 , n369 ); 
nor ( n640 , n16 , n207 ); 
not ( n641 , n640 ); 
nand ( n642 , n357 , n641 ); 
nand ( n643 , n639 , n642 ); 
not ( n644 , n641 ); 
nand ( n645 , n644 , n642 ); 
not ( n646 , n640 ); 
not ( n647 , n357 ); 
nor ( n648 , n647 , n640 ); 
nand ( n649 , n646 , n369 , n648 ); 
nand ( n650 , n643 , n645 , n649 ); 
and ( n651 , n278 , n650 ); 
nand ( n652 , n584 , n612 , n638 , n651 ); 
nor ( n653 , n547 , n652 ); 
not ( n654 , n163 ); 
not ( n655 , n79 ); 
nand ( n656 , n655 , n578 ); 
not ( n657 , n573 ); 
nand ( n658 , n657 , n79 , n574 ); 
nand ( n659 , n656 , n579 , n658 ); 
not ( n660 , n91 ); 
nand ( n661 , n660 , n564 ); 
not ( n662 , n562 ); 
nand ( n663 , n662 , n91 , n563 ); 
nand ( n664 , n661 , n568 , n663 ); 
or ( n665 , n43 , n551 ); 
not ( n666 , n550 ); 
nand ( n667 , n666 , n43 , n551 ); 
nand ( n668 , n665 , n556 , n667 ); 
nand ( n669 , n659 , n664 , n668 ); 
not ( n670 , n669 ); 
not ( n671 , n55 ); 
nand ( n672 , n671 , n601 ); 
not ( n673 , n606 ); 
nand ( n674 , n673 , n55 , n608 ); 
nand ( n675 , n672 , n605 , n674 ); 
nand ( n676 , n159 , n675 ); 
not ( n677 , n676 ); 
not ( n678 , n1 ); 
nand ( n679 , n678 , n616 ); 
not ( n680 , n621 ); 
nand ( n681 , n680 , n1 , n623 ); 
nand ( n682 , n679 , n620 , n681 ); 
not ( n683 , n358 ); 
nand ( n684 , n683 , n642 ); 
not ( n685 , n640 ); 
nand ( n686 , n685 , n358 , n648 ); 
nand ( n687 , n684 , n645 , n686 ); 
and ( n688 , n682 , n687 ); 
not ( n689 , n67 ); 
nand ( n690 , n689 , n588 ); 
not ( n691 , n594 ); 
not ( n692 , n588 ); 
nand ( n693 , n691 , n67 , n692 ); 
nand ( n694 , n690 , n592 , n693 ); 
not ( n695 , n355 ); 
nand ( n696 , n695 , n629 ); 
not ( n697 , n627 ); 
nand ( n698 , n697 , n355 , n635 ); 
nand ( n699 , n696 , n632 , n698 ); 
nand ( n700 , n694 , n699 ); 
not ( n701 , n700 ); 
nand ( n702 , n670 , n677 , n688 , n701 ); 
nor ( n703 , n654 , n702 ); 
or ( n704 , n653 , n703 ); 
and ( n705 , n349 , n544 ); 
nand ( n706 , n704 , n705 ); 
nand ( n707 , n546 , n706 ); 
not ( n708 , n345 ); 
not ( n709 , n362 ); 
nor ( n710 , n709 , n16 ); 
nand ( n711 , n708 , n710 ); 
not ( n712 , n710 ); 
not ( n713 , n712 ); 
not ( n714 , n16 ); 
nand ( n715 , n714 , n366 ); 
not ( n716 , n16 ); 
nand ( n717 , n716 , n365 ); 
not ( n718 , n717 ); 
not ( n719 , n364 ); 
nor ( n720 , n719 , n16 ); 
not ( n721 , n16 ); 
nand ( n722 , n721 , n363 ); 
not ( n723 , n722 ); 
not ( n724 , n16 ); 
nand ( n725 , n724 , n361 ); 
not ( n726 , n344 ); 
nor ( n727 , n726 , n16 ); 
not ( n728 , n360 ); 
nor ( n729 , n728 , n16 ); 
nand ( n730 , n727 , n729 ); 
nor ( n731 , n725 , n730 ); 
and ( n732 , n720 , n723 , n731 ); 
nand ( n733 , n718 , n732 ); 
nor ( n734 , n715 , n733 ); 
not ( n735 , n734 ); 
not ( n736 , n735 ); 
or ( n737 , n713 , n736 ); 
not ( n738 , n710 ); 
not ( n739 , n734 ); 
or ( n740 , n738 , n739 ); 
nand ( n741 , n740 , n345 ); 
not ( n742 , n741 ); 
nand ( n743 , n737 , n742 ); 
and ( n744 , n711 , n743 ); 
not ( n745 , n16 ); 
nand ( n746 , n745 , n346 ); 
not ( n747 , n746 ); 
nor ( n748 , n744 , n747 ); 
not ( n749 , n91 ); 
not ( n750 , n6 ); 
xor ( n751 , n2 , n3 ); 
not ( n752 , n751 ); 
and ( n753 , n750 , n5 , n4 , n752 ); 
buf ( n754 , n753 ); 
not ( n755 , n754 ); 
or ( n756 , n749 , n755 ); 
and ( n757 , n6 , n5 , n4 , n752 ); 
buf ( n758 , n757 ); 
nand ( n759 , n92 , n758 ); 
nand ( n760 , n756 , n759 ); 
nor ( n761 , n4 , n751 ); 
and ( n762 , n6 , n5 , n761 ); 
buf ( n763 , n762 ); 
nand ( n764 , n93 , n763 ); 
and ( n765 , n750 , n5 , n761 ); 
buf ( n766 , n765 ); 
nand ( n767 , n95 , n766 ); 
not ( n768 , n5 ); 
not ( n769 , n4 ); 
nand ( n770 , n6 , n768 , n769 , n752 ); 
not ( n771 , n770 ); 
nand ( n772 , n94 , n771 ); 
nand ( n773 , n764 , n767 , n772 ); 
nor ( n774 , n760 , n773 ); 
not ( n775 , n12 ); 
nor ( n776 , n11 , n13 ); 
and ( n777 , n775 , n776 ); 
buf ( n778 , n777 ); 
or ( n779 , n774 , n778 ); 
buf ( n780 , n777 ); 
not ( n781 , n17 ); 
nor ( n782 , n781 , n16 ); 
not ( n783 , n782 ); 
not ( n784 , n16 ); 
nand ( n785 , n784 , n15 ); 
nand ( n786 , n783 , n785 ); 
not ( n787 , n786 ); 
nand ( n788 , n98 , n787 ); 
not ( n789 , n782 ); 
buf ( n790 , n789 ); 
not ( n791 , n790 ); 
nand ( n792 , n97 , n791 ); 
not ( n793 , n782 ); 
not ( n794 , n785 ); 
nand ( n795 , n793 , n794 ); 
not ( n796 , n795 ); 
nand ( n797 , n96 , n796 ); 
and ( n798 , n788 , n792 , n797 ); 
nor ( n799 , n20 , n21 ); 
or ( n800 , n16 , n799 ); 
buf ( n801 , n800 ); 
nor ( n802 , n798 , n801 ); 
not ( n803 , n802 ); 
not ( n804 , n99 ); 
not ( n805 , n16 ); 
nand ( n806 , n805 , n25 ); 
not ( n807 , n16 ); 
nand ( n808 , n807 , n26 ); 
nand ( n809 , n806 , n808 ); 
not ( n810 , n23 ); 
nor ( n811 , n810 , n16 ); 
not ( n812 , n811 ); 
not ( n813 , n16 ); 
not ( n814 , n24 ); 
nand ( n815 , n813 , n814 ); 
nand ( n816 , n812 , n815 ); 
nor ( n817 , n809 , n816 ); 
buf ( n818 , n817 ); 
not ( n819 , n818 ); 
or ( n820 , n804 , n819 ); 
nor ( n821 , n16 , n24 ); 
nand ( n822 , n806 , n808 , n811 , n821 ); 
not ( n823 , n822 ); 
buf ( n824 , n823 ); 
nand ( n825 , n101 , n824 ); 
nand ( n826 , n820 , n825 ); 
not ( n827 , n100 ); 
not ( n828 , n808 ); 
nand ( n829 , n828 , n806 ); 
not ( n830 , n16 ); 
nand ( n831 , n830 , n23 ); 
nand ( n832 , n831 , n821 ); 
nor ( n833 , n829 , n832 ); 
buf ( n834 , n833 ); 
not ( n835 , n834 ); 
or ( n836 , n827 , n835 ); 
not ( n837 , n806 ); 
nand ( n838 , n837 , n808 ); 
nand ( n839 , n831 , n821 ); 
nor ( n840 , n838 , n839 ); 
buf ( n841 , n840 ); 
nand ( n842 , n102 , n841 ); 
nand ( n843 , n836 , n842 ); 
or ( n844 , n826 , n843 ); 
not ( n845 , n801 ); 
not ( n846 , n845 ); 
nand ( n847 , n844 , n846 ); 
nand ( n848 , n803 , n847 ); 
nand ( n849 , n780 , n848 ); 
nand ( n850 , n779 , n849 ); 
not ( n851 , n47 ); 
buf ( n852 , n765 ); 
not ( n853 , n852 ); 
or ( n854 , n851 , n853 ); 
nand ( n855 , n46 , n771 ); 
nand ( n856 , n854 , n855 ); 
nand ( n857 , n45 , n763 ); 
nand ( n858 , n44 , n758 ); 
nand ( n859 , n43 , n754 ); 
nand ( n860 , n857 , n858 , n859 ); 
nor ( n861 , n856 , n860 ); 
or ( n862 , n778 , n861 ); 
nand ( n863 , n49 , n791 ); 
nand ( n864 , n50 , n787 ); 
nand ( n865 , n48 , n796 ); 
and ( n866 , n863 , n864 , n865 ); 
nor ( n867 , n866 , n801 ); 
not ( n868 , n867 ); 
not ( n869 , n51 ); 
not ( n870 , n818 ); 
or ( n871 , n869 , n870 ); 
nand ( n872 , n52 , n841 ); 
nand ( n873 , n871 , n872 ); 
not ( n874 , n53 ); 
not ( n875 , n834 ); 
or ( n876 , n874 , n875 ); 
buf ( n877 , n823 ); 
nand ( n878 , n54 , n877 ); 
nand ( n879 , n876 , n878 ); 
or ( n880 , n873 , n879 ); 
nand ( n881 , n880 , n846 ); 
nand ( n882 , n868 , n881 ); 
nand ( n883 , n778 , n882 ); 
nand ( n884 , n862 , n883 ); 
not ( n885 , n59 ); 
not ( n886 , n852 ); 
or ( n887 , n885 , n886 ); 
nand ( n888 , n58 , n771 ); 
nand ( n889 , n887 , n888 ); 
nand ( n890 , n57 , n763 ); 
nand ( n891 , n56 , n758 ); 
nand ( n892 , n55 , n754 ); 
nand ( n893 , n890 , n891 , n892 ); 
nor ( n894 , n889 , n893 ); 
or ( n895 , n778 , n894 ); 
nand ( n896 , n62 , n787 ); 
nand ( n897 , n61 , n791 ); 
nand ( n898 , n60 , n796 ); 
and ( n899 , n896 , n897 , n898 ); 
nor ( n900 , n899 , n801 ); 
not ( n901 , n900 ); 
not ( n902 , n63 ); 
not ( n903 , n818 ); 
or ( n904 , n902 , n903 ); 
nand ( n905 , n65 , n824 ); 
nand ( n906 , n904 , n905 ); 
not ( n907 , n64 ); 
not ( n908 , n834 ); 
or ( n909 , n907 , n908 ); 
nand ( n910 , n66 , n841 ); 
nand ( n911 , n909 , n910 ); 
or ( n912 , n906 , n911 ); 
buf ( n913 , n801 ); 
nand ( n914 , n912 , n913 ); 
nand ( n915 , n901 , n914 ); 
nand ( n916 , n778 , n915 ); 
nand ( n917 , n895 , n916 ); 
not ( n918 , n71 ); 
not ( n919 , n852 ); 
or ( n920 , n918 , n919 ); 
nand ( n921 , n70 , n771 ); 
nand ( n922 , n920 , n921 ); 
nand ( n923 , n69 , n763 ); 
nand ( n924 , n68 , n758 ); 
nand ( n925 , n67 , n754 ); 
nand ( n926 , n923 , n924 , n925 ); 
nor ( n927 , n922 , n926 ); 
or ( n928 , n778 , n927 ); 
nand ( n929 , n74 , n787 ); 
nand ( n930 , n73 , n791 ); 
nand ( n931 , n72 , n796 ); 
and ( n932 , n929 , n930 , n931 ); 
nor ( n933 , n932 , n801 ); 
not ( n934 , n933 ); 
not ( n935 , n77 ); 
not ( n936 , n834 ); 
or ( n937 , n935 , n936 ); 
nand ( n938 , n75 , n818 ); 
nand ( n939 , n937 , n938 ); 
not ( n940 , n78 ); 
and ( n941 , n837 , n808 , n831 , n821 ); 
buf ( n942 , n941 ); 
not ( n943 , n942 ); 
or ( n944 , n940 , n943 ); 
nand ( n945 , n76 , n877 ); 
nand ( n946 , n944 , n945 ); 
or ( n947 , n939 , n946 ); 
nand ( n948 , n947 , n913 ); 
nand ( n949 , n934 , n948 ); 
nand ( n950 , n778 , n949 ); 
nand ( n951 , n928 , n950 ); 
not ( n952 , n83 ); 
not ( n953 , n852 ); 
or ( n954 , n952 , n953 ); 
nand ( n955 , n82 , n771 ); 
nand ( n956 , n954 , n955 ); 
nand ( n957 , n81 , n763 ); 
nand ( n958 , n80 , n758 ); 
nand ( n959 , n79 , n754 ); 
nand ( n960 , n957 , n958 , n959 ); 
nor ( n961 , n956 , n960 ); 
or ( n962 , n778 , n961 ); 
nand ( n963 , n85 , n791 ); 
nand ( n964 , n86 , n787 ); 
nand ( n965 , n84 , n796 ); 
and ( n966 , n963 , n964 , n965 ); 
nor ( n967 , n966 , n801 ); 
not ( n968 , n967 ); 
not ( n969 , n87 ); 
not ( n970 , n818 ); 
or ( n971 , n969 , n970 ); 
nand ( n972 , n90 , n841 ); 
nand ( n973 , n971 , n972 ); 
not ( n974 , n88 ); 
not ( n975 , n834 ); 
or ( n976 , n974 , n975 ); 
nand ( n977 , n89 , n877 ); 
nand ( n978 , n976 , n977 ); 
or ( n979 , n973 , n978 ); 
nand ( n980 , n979 , n913 ); 
nand ( n981 , n968 , n980 ); 
nand ( n982 , n778 , n981 ); 
nand ( n983 , n962 , n982 ); 
and ( n984 , n8 , n763 ); 
not ( n985 , n1 ); 
not ( n986 , n754 ); 
or ( n987 , n985 , n986 ); 
nand ( n988 , n7 , n758 ); 
nand ( n989 , n987 , n988 ); 
not ( n990 , n10 ); 
not ( n991 , n852 ); 
or ( n992 , n990 , n991 ); 
nand ( n993 , n9 , n771 ); 
nand ( n994 , n992 , n993 ); 
nor ( n995 , n984 , n989 , n994 ); 
or ( n996 , n995 , n778 ); 
buf ( n997 , n801 ); 
not ( n998 , n997 ); 
not ( n999 , n29 ); 
not ( n1000 , n942 ); 
or ( n1001 , n999 , n1000 ); 
nand ( n1002 , n30 , n877 ); 
nand ( n1003 , n1001 , n1002 ); 
nor ( n1004 , n809 , n816 ); 
not ( n1005 , n1004 ); 
not ( n1006 , n28 ); 
nor ( n1007 , n1005 , n1006 ); 
not ( n1008 , n1007 ); 
and ( n1009 , n806 , n828 , n831 , n821 ); 
nand ( n1010 , n27 , n1009 ); 
not ( n1011 , n1010 ); 
or ( n1012 , n1008 , n1011 ); 
or ( n1013 , n1007 , n1010 ); 
nand ( n1014 , n1012 , n1013 ); 
nor ( n1015 , n1003 , n1014 ); 
or ( n1016 , n998 , n1015 ); 
not ( n1017 , n789 ); 
nand ( n1018 , n18 , n1017 ); 
not ( n1019 , n1018 ); 
not ( n1020 , n786 ); 
nand ( n1021 , n19 , n1020 ); 
not ( n1022 , n1021 ); 
or ( n1023 , n1019 , n1022 ); 
and ( n1024 , n14 , n796 ); 
nor ( n1025 , 1'b0 , n1024 ); 
nand ( n1026 , n1023 , n1025 ); 
nand ( n1027 , n845 , n1026 ); 
nand ( n1028 , n1016 , n1027 ); 
nand ( n1029 , n778 , n1028 ); 
nand ( n1030 , n996 , n1029 ); 
not ( n1031 , n106 ); 
not ( n1032 , n771 ); 
or ( n1033 , n1031 , n1032 ); 
nand ( n1034 , n105 , n763 ); 
nand ( n1035 , n1033 , n1034 ); 
not ( n1036 , n103 ); 
not ( n1037 , n754 ); 
or ( n1038 , n1036 , n1037 ); 
nand ( n1039 , n104 , n758 ); 
nand ( n1040 , n1038 , n1039 ); 
not ( n1041 , n108 ); 
not ( n1042 , n766 ); 
or ( n1043 , n1041 , n1042 ); 
not ( n1044 , n16 ); 
not ( n1045 , n751 ); 
nand ( n1046 , n1045 , n750 , n768 , n769 ); 
not ( n1047 , n1046 ); 
nand ( n1048 , n107 , n1044 , n1047 ); 
nand ( n1049 , n1043 , n1048 ); 
nor ( n1050 , n1035 , n1040 , n1049 ); 
or ( n1051 , n1050 , n778 ); 
not ( n1052 , n786 ); 
and ( n1053 , n84 , n1052 ); 
not ( n1054 , n110 ); 
not ( n1055 , n796 ); 
or ( n1056 , n1054 , n1055 ); 
not ( n1057 , n789 ); 
nand ( n1058 , n109 , n1057 ); 
nand ( n1059 , n1056 , n1058 ); 
nor ( n1060 , n1053 , n1059 ); 
nor ( n1061 , n801 , n1060 ); 
not ( n1062 , n1061 ); 
not ( n1063 , n111 ); 
not ( n1064 , n818 ); 
or ( n1065 , n1063 , n1064 ); 
nand ( n1066 , n113 , n824 ); 
nand ( n1067 , n1065 , n1066 ); 
not ( n1068 , n112 ); 
not ( n1069 , n834 ); 
or ( n1070 , n1068 , n1069 ); 
nand ( n1071 , n114 , n841 ); 
nand ( n1072 , n1070 , n1071 ); 
or ( n1073 , n1067 , n1072 ); 
not ( n1074 , n845 ); 
nand ( n1075 , n1073 , n1074 ); 
nand ( n1076 , n1062 , n1075 ); 
nand ( n1077 , n780 , n1076 ); 
nand ( n1078 , n1051 , n1077 ); 
not ( n1079 , n118 ); 
not ( n1080 , n771 ); 
or ( n1081 , n1079 , n1080 ); 
nand ( n1082 , n117 , n763 ); 
nand ( n1083 , n1081 , n1082 ); 
not ( n1084 , n115 ); 
not ( n1085 , n754 ); 
or ( n1086 , n1084 , n1085 ); 
nand ( n1087 , n116 , n758 ); 
nand ( n1088 , n1086 , n1087 ); 
not ( n1089 , n120 ); 
not ( n1090 , n852 ); 
or ( n1091 , n1089 , n1090 ); 
nand ( n1092 , n119 , n1044 , n1047 ); 
nand ( n1093 , n1091 , n1092 ); 
nor ( n1094 , n1083 , n1088 , n1093 ); 
or ( n1095 , n1094 , n778 ); 
and ( n1096 , n123 , n1052 ); 
not ( n1097 , n121 ); 
not ( n1098 , n796 ); 
or ( n1099 , n1097 , n1098 ); 
nand ( n1100 , n122 , n1057 ); 
nand ( n1101 , n1099 , n1100 ); 
nor ( n1102 , n1096 , n1101 ); 
nor ( n1103 , n801 , n1102 ); 
not ( n1104 , n1103 ); 
not ( n1105 , n124 ); 
not ( n1106 , n818 ); 
or ( n1107 , n1105 , n1106 ); 
nand ( n1108 , n127 , n824 ); 
nand ( n1109 , n1107 , n1108 ); 
not ( n1110 , n126 ); 
not ( n1111 , n834 ); 
or ( n1112 , n1110 , n1111 ); 
nand ( n1113 , n125 , n841 ); 
nand ( n1114 , n1112 , n1113 ); 
or ( n1115 , n1109 , n1114 ); 
buf ( n1116 , n801 ); 
nand ( n1117 , n1115 , n1116 ); 
nand ( n1118 , n1104 , n1117 ); 
nand ( n1119 , n780 , n1118 ); 
nand ( n1120 , n1095 , n1119 ); 
nand ( n1121 , n131 , n763 ); 
nand ( n1122 , n133 , n758 ); 
nand ( n1123 , n132 , n754 ); 
nand ( n1124 , n1121 , n1122 , n1123 ); 
nand ( n1125 , n130 , n1044 , n1047 ); 
nand ( n1126 , n129 , n766 ); 
nand ( n1127 , n128 , n771 ); 
nand ( n1128 , n1125 , n1126 , n1127 ); 
nor ( n1129 , n1124 , n1128 ); 
or ( n1130 , n1129 , n778 ); 
nand ( n1131 , n60 , n787 ); 
nand ( n1132 , n134 , n791 ); 
nand ( n1133 , n135 , n796 ); 
and ( n1134 , n1131 , n1132 , n1133 ); 
nor ( n1135 , n1134 , n801 ); 
not ( n1136 , n1135 ); 
not ( n1137 , n136 ); 
not ( n1138 , n818 ); 
or ( n1139 , n1137 , n1138 ); 
nand ( n1140 , n138 , n824 ); 
nand ( n1141 , n1139 , n1140 ); 
not ( n1142 , n137 ); 
not ( n1143 , n834 ); 
or ( n1144 , n1142 , n1143 ); 
nand ( n1145 , n139 , n841 ); 
nand ( n1146 , n1144 , n1145 ); 
or ( n1147 , n1141 , n1146 ); 
nand ( n1148 , n1147 , n913 ); 
nand ( n1149 , n1136 , n1148 ); 
nand ( n1150 , n778 , n1149 ); 
nand ( n1151 , n1130 , n1150 ); 
not ( n1152 , n144 ); 
not ( n1153 , n852 ); 
or ( n1154 , n1152 , n1153 ); 
nand ( n1155 , n143 , n771 ); 
nand ( n1156 , n1154 , n1155 ); 
nand ( n1157 , n142 , n763 ); 
nand ( n1158 , n141 , n758 ); 
nand ( n1159 , n140 , n754 ); 
nand ( n1160 , n1157 , n1158 , n1159 ); 
nor ( n1161 , n1156 , n1160 ); 
or ( n1162 , n778 , n1161 ); 
not ( n1163 , n790 ); 
nand ( n1164 , n38 , n1163 ); 
nand ( n1165 , n795 , n786 ); 
buf ( n1166 , n1165 ); 
nand ( n1167 , n145 , n1166 ); 
and ( n1168 , n1164 , n1167 ); 
nor ( n1169 , n1168 , n801 ); 
not ( n1170 , n1169 ); 
not ( n1171 , n146 ); 
not ( n1172 , n818 ); 
or ( n1173 , n1171 , n1172 ); 
nand ( n1174 , n148 , n824 ); 
nand ( n1175 , n1173 , n1174 ); 
not ( n1176 , n147 ); 
not ( n1177 , n834 ); 
or ( n1178 , n1176 , n1177 ); 
nand ( n1179 , n149 , n841 ); 
nand ( n1180 , n1178 , n1179 ); 
or ( n1181 , n1175 , n1180 ); 
nand ( n1182 , n1181 , n913 ); 
nand ( n1183 , n1170 , n1182 ); 
nand ( n1184 , n778 , n1183 ); 
nand ( n1185 , n1162 , n1184 ); 
not ( n1186 , n165 ); 
not ( n1187 , n771 ); 
or ( n1188 , n1186 , n1187 ); 
and ( n1189 , n166 , n1044 , n1047 ); 
not ( n1190 , n16 ); 
not ( n1191 , n167 ); 
and ( n1192 , n1190 , n1191 ); 
not ( n1193 , n751 ); 
nor ( n1194 , n5 , n6 ); 
nand ( n1195 , n1193 , n1194 , n4 ); 
nor ( n1196 , n1192 , n1195 ); 
nor ( n1197 , n1189 , n1196 ); 
nand ( n1198 , n1188 , n1197 ); 
not ( n1199 , n163 ); 
not ( n1200 , n754 ); 
or ( n1201 , n1199 , n1200 ); 
nand ( n1202 , n164 , n758 ); 
nand ( n1203 , n1201 , n1202 ); 
not ( n1204 , n161 ); 
not ( n1205 , n852 ); 
or ( n1206 , n1204 , n1205 ); 
nand ( n1207 , n162 , n763 ); 
nand ( n1208 , n1206 , n1207 ); 
nor ( n1209 , n1198 , n1203 , n1208 ); 
or ( n1210 , n1209 , n778 ); 
buf ( n1211 , n1057 ); 
nand ( n1212 , n121 , n1211 ); 
nand ( n1213 , n168 , n1166 ); 
and ( n1214 , n1212 , n1213 ); 
nor ( n1215 , n1214 , n801 ); 
not ( n1216 , n1215 ); 
not ( n1217 , n170 ); 
not ( n1218 , n834 ); 
or ( n1219 , n1217 , n1218 ); 
nand ( n1220 , n172 , n942 ); 
nand ( n1221 , n1219 , n1220 ); 
not ( n1222 , n169 ); 
not ( n1223 , n818 ); 
or ( n1224 , n1222 , n1223 ); 
nand ( n1225 , n171 , n824 ); 
nand ( n1226 , n1224 , n1225 ); 
or ( n1227 , n1221 , n1226 ); 
nand ( n1228 , n1227 , n997 ); 
nand ( n1229 , n1216 , n1228 ); 
nand ( n1230 , n778 , n1229 ); 
nand ( n1231 , n1210 , n1230 ); 
nand ( n1232 , n246 , n1044 , n1047 ); 
nand ( n1233 , n244 , n771 ); 
not ( n1234 , n1195 ); 
nand ( n1235 , n566 , n1234 ); 
nand ( n1236 , n1232 , n1233 , n1235 ); 
not ( n1237 , n249 ); 
not ( n1238 , n754 ); 
or ( n1239 , n1237 , n1238 ); 
nand ( n1240 , n250 , n758 ); 
nand ( n1241 , n1239 , n1240 ); 
not ( n1242 , n247 ); 
not ( n1243 , n766 ); 
or ( n1244 , n1242 , n1243 ); 
nand ( n1245 , n248 , n763 ); 
nand ( n1246 , n1244 , n1245 ); 
nor ( n1247 , n1236 , n1241 , n1246 ); 
or ( n1248 , n1247 , n778 ); 
nand ( n1249 , n96 , n1211 ); 
nand ( n1250 , n251 , n1166 ); 
and ( n1251 , n1249 , n1250 ); 
nor ( n1252 , n1251 , n801 ); 
not ( n1253 , n1252 ); 
not ( n1254 , n252 ); 
not ( n1255 , n818 ); 
or ( n1256 , n1254 , n1255 ); 
nand ( n1257 , n255 , n942 ); 
nand ( n1258 , n1256 , n1257 ); 
not ( n1259 , n253 ); 
not ( n1260 , n834 ); 
or ( n1261 , n1259 , n1260 ); 
nand ( n1262 , n254 , n877 ); 
nand ( n1263 , n1261 , n1262 ); 
or ( n1264 , n1258 , n1263 ); 
nand ( n1265 , n1264 , n1116 ); 
nand ( n1266 , n1253 , n1265 ); 
nand ( n1267 , n780 , n1266 ); 
nand ( n1268 , n1248 , n1267 ); 
not ( n1269 , n187 ); 
not ( n1270 , n852 ); 
or ( n1271 , n1269 , n1270 ); 
nand ( n1272 , n186 , n771 ); 
nand ( n1273 , n1271 , n1272 ); 
nand ( n1274 , n185 , n763 ); 
nand ( n1275 , n184 , n758 ); 
nand ( n1276 , n183 , n754 ); 
nand ( n1277 , n1274 , n1275 , n1276 ); 
nor ( n1278 , n1273 , n1277 ); 
or ( n1279 , n778 , n1278 ); 
nand ( n1280 , n188 , n1163 ); 
nand ( n1281 , n189 , n1166 ); 
and ( n1282 , n1280 , n1281 ); 
nor ( n1283 , n1282 , n801 ); 
not ( n1284 , n1283 ); 
not ( n1285 , n191 ); 
not ( n1286 , n834 ); 
or ( n1287 , n1285 , n1286 ); 
nand ( n1288 , n190 , n818 ); 
nand ( n1289 , n1287 , n1288 ); 
not ( n1290 , n193 ); 
not ( n1291 , n942 ); 
or ( n1292 , n1290 , n1291 ); 
nand ( n1293 , n192 , n877 ); 
nand ( n1294 , n1292 , n1293 ); 
or ( n1295 , n1289 , n1294 ); 
nand ( n1296 , n1295 , n846 ); 
nand ( n1297 , n1284 , n1296 ); 
nand ( n1298 , n780 , n1297 ); 
nand ( n1299 , n1279 , n1298 ); 
nand ( n1300 , n281 , n771 ); 
nand ( n1301 , n280 , n758 ); 
nand ( n1302 , n159 , n754 ); 
nand ( n1303 , n1300 , n1301 , n1302 ); 
not ( n1304 , n627 ); 
not ( n1305 , n1195 ); 
and ( n1306 , n1304 , n1305 ); 
and ( n1307 , n282 , n1047 ); 
nor ( n1308 , n1306 , n1307 ); 
nand ( n1309 , n279 , n763 ); 
nand ( n1310 , n278 , n766 ); 
nand ( n1311 , n1308 , n1309 , n1310 ); 
nor ( n1312 , n1303 , n1311 ); 
or ( n1313 , n1312 , n778 ); 
nand ( n1314 , n123 , n1211 ); 
nand ( n1315 , n284 , n1166 ); 
and ( n1316 , n1314 , n1315 ); 
nor ( n1317 , n1316 , n801 ); 
not ( n1318 , n1317 ); 
not ( n1319 , n287 ); 
not ( n1320 , n834 ); 
or ( n1321 , n1319 , n1320 ); 
nand ( n1322 , n286 , n942 ); 
nand ( n1323 , n1321 , n1322 ); 
not ( n1324 , n285 ); 
not ( n1325 , n818 ); 
or ( n1326 , n1324 , n1325 ); 
nand ( n1327 , n288 , n824 ); 
nand ( n1328 , n1326 , n1327 ); 
or ( n1329 , n1323 , n1328 ); 
nand ( n1330 , n1329 , n997 ); 
nand ( n1331 , n1318 , n1330 ); 
nand ( n1332 , n778 , n1331 ); 
nand ( n1333 , n1313 , n1332 ); 
nand ( n1334 , n304 , n771 ); 
nand ( n1335 , n303 , n758 ); 
nand ( n1336 , n302 , n754 ); 
nand ( n1337 , n1334 , n1335 , n1336 ); 
not ( n1338 , n606 ); 
not ( n1339 , n1195 ); 
and ( n1340 , n1338 , n1339 ); 
and ( n1341 , n305 , n1047 ); 
nor ( n1342 , n1340 , n1341 ); 
nand ( n1343 , n301 , n763 ); 
nand ( n1344 , n300 , n766 ); 
nand ( n1345 , n1342 , n1343 , n1344 ); 
nor ( n1346 , n1337 , n1345 ); 
or ( n1347 , n1346 , n778 ); 
nand ( n1348 , n307 , n1166 ); 
nand ( n1349 , n60 , n1163 ); 
and ( n1350 , n1348 , n1349 ); 
nor ( n1351 , n1350 , n801 ); 
not ( n1352 , n1351 ); 
not ( n1353 , n311 ); 
not ( n1354 , n834 ); 
or ( n1355 , n1353 , n1354 ); 
nand ( n1356 , n310 , n818 ); 
nand ( n1357 , n1355 , n1356 ); 
not ( n1358 , n309 ); 
not ( n1359 , n942 ); 
or ( n1360 , n1358 , n1359 ); 
nand ( n1361 , n308 , n877 ); 
nand ( n1362 , n1360 , n1361 ); 
or ( n1363 , n1357 , n1362 ); 
nand ( n1364 , n1363 , n1074 ); 
nand ( n1365 , n1352 , n1364 ); 
nand ( n1366 , n780 , n1365 ); 
nand ( n1367 , n1347 , n1366 ); 
nand ( n1368 , n316 , n1044 , n1047 ); 
nand ( n1369 , n317 , n771 ); 
nand ( n1370 , n576 , n1234 ); 
nand ( n1371 , n1368 , n1369 , n1370 ); 
not ( n1372 , n314 ); 
not ( n1373 , n754 ); 
or ( n1374 , n1372 , n1373 ); 
nand ( n1375 , n315 , n758 ); 
nand ( n1376 , n1374 , n1375 ); 
not ( n1377 , n312 ); 
not ( n1378 , n766 ); 
or ( n1379 , n1377 , n1378 ); 
nand ( n1380 , n313 , n763 ); 
nand ( n1381 , n1379 , n1380 ); 
nor ( n1382 , n1371 , n1376 , n1381 ); 
or ( n1383 , n1382 , n778 ); 
nand ( n1384 , n84 , n1211 ); 
nand ( n1385 , n319 , n1166 ); 
and ( n1386 , n1384 , n1385 ); 
nor ( n1387 , n1386 , n801 ); 
not ( n1388 , n1387 ); 
not ( n1389 , n320 ); 
not ( n1390 , n818 ); 
or ( n1391 , n1389 , n1390 ); 
nand ( n1392 , n322 , n824 ); 
nand ( n1393 , n1391 , n1392 ); 
not ( n1394 , n321 ); 
not ( n1395 , n834 ); 
or ( n1396 , n1394 , n1395 ); 
nand ( n1397 , n323 , n841 ); 
nand ( n1398 , n1396 , n1397 ); 
or ( n1399 , n1393 , n1398 ); 
nand ( n1400 , n1399 , n1074 ); 
nand ( n1401 , n1388 , n1400 ); 
nand ( n1402 , n780 , n1401 ); 
nand ( n1403 , n1383 , n1402 ); 
not ( n1404 , n328 ); 
not ( n1405 , n771 ); 
or ( n1406 , n1404 , n1405 ); 
and ( n1407 , n329 , n1044 , n1047 ); 
not ( n1408 , n16 ); 
not ( n1409 , n330 ); 
and ( n1410 , n1408 , n1409 ); 
nor ( n1411 , n1410 , n1195 ); 
nor ( n1412 , n1407 , n1411 ); 
nand ( n1413 , n1406 , n1412 ); 
not ( n1414 , n326 ); 
not ( n1415 , n754 ); 
or ( n1416 , n1414 , n1415 ); 
nand ( n1417 , n327 , n758 ); 
nand ( n1418 , n1416 , n1417 ); 
not ( n1419 , n324 ); 
not ( n1420 , n766 ); 
or ( n1421 , n1419 , n1420 ); 
nand ( n1422 , n325 , n763 ); 
nand ( n1423 , n1421 , n1422 ); 
nor ( n1424 , n1413 , n1418 , n1423 ); 
or ( n1425 , n1424 , n778 ); 
nand ( n1426 , n331 , n1166 ); 
nand ( n1427 , n110 , n1211 ); 
and ( n1428 , n1426 , n1427 ); 
nor ( n1429 , n1428 , n801 ); 
not ( n1430 , n1429 ); 
not ( n1431 , n333 ); 
not ( n1432 , n834 ); 
or ( n1433 , n1431 , n1432 ); 
nand ( n1434 , n335 , n942 ); 
nand ( n1435 , n1433 , n1434 ); 
not ( n1436 , n332 ); 
not ( n1437 , n818 ); 
or ( n1438 , n1436 , n1437 ); 
nand ( n1439 , n334 , n824 ); 
nand ( n1440 , n1438 , n1439 ); 
or ( n1441 , n1435 , n1440 ); 
nand ( n1442 , n1441 , n1116 ); 
nand ( n1443 , n1430 , n1442 ); 
nand ( n1444 , n778 , n1443 ); 
nand ( n1445 , n1425 , n1444 ); 
and ( n1446 , n175 , n763 ); 
not ( n1447 , n173 ); 
not ( n1448 , n754 ); 
or ( n1449 , n1447 , n1448 ); 
nand ( n1450 , n174 , n758 ); 
nand ( n1451 , n1449 , n1450 ); 
not ( n1452 , n177 ); 
not ( n1453 , n766 ); 
or ( n1454 , n1452 , n1453 ); 
nand ( n1455 , n176 , n771 ); 
nand ( n1456 , n1454 , n1455 ); 
nor ( n1457 , n1446 , n1451 , n1456 ); 
or ( n1458 , n1457 , n778 ); 
nand ( n1459 , n135 , n1163 ); 
nand ( n1460 , n178 , n1166 ); 
and ( n1461 , n1459 , n1460 ); 
nor ( n1462 , n1461 , n801 ); 
not ( n1463 , n1462 ); 
not ( n1464 , n179 ); 
not ( n1465 , n818 ); 
or ( n1466 , n1464 , n1465 ); 
nand ( n1467 , n182 , n841 ); 
nand ( n1468 , n1466 , n1467 ); 
not ( n1469 , n180 ); 
not ( n1470 , n834 ); 
or ( n1471 , n1469 , n1470 ); 
nand ( n1472 , n181 , n877 ); 
nand ( n1473 , n1471 , n1472 ); 
or ( n1474 , n1468 , n1473 ); 
nand ( n1475 , n1474 , n913 ); 
nand ( n1476 , n1463 , n1475 ); 
nand ( n1477 , n780 , n1476 ); 
nand ( n1478 , n1458 , n1477 ); 
and ( n1479 , n269 , n763 ); 
not ( n1480 , n267 ); 
not ( n1481 , n754 ); 
or ( n1482 , n1480 , n1481 ); 
nand ( n1483 , n268 , n758 ); 
nand ( n1484 , n1482 , n1483 ); 
not ( n1485 , n271 ); 
not ( n1486 , n766 ); 
or ( n1487 , n1485 , n1486 ); 
nand ( n1488 , n270 , n771 ); 
nand ( n1489 , n1487 , n1488 ); 
nor ( n1490 , n1479 , n1484 , n1489 ); 
or ( n1491 , n1490 , n778 ); 
nand ( n1492 , n272 , n1163 ); 
nand ( n1493 , n273 , n1166 ); 
and ( n1494 , n1492 , n1493 ); 
nor ( n1495 , n1494 , n801 ); 
not ( n1496 , n1495 ); 
not ( n1497 , n274 ); 
not ( n1498 , n818 ); 
or ( n1499 , n1497 , n1498 ); 
nand ( n1500 , n277 , n841 ); 
nand ( n1501 , n1499 , n1500 ); 
not ( n1502 , n275 ); 
not ( n1503 , n834 ); 
or ( n1504 , n1502 , n1503 ); 
nand ( n1505 , n276 , n877 ); 
nand ( n1506 , n1504 , n1505 ); 
or ( n1507 , n1501 , n1506 ); 
nand ( n1508 , n1507 , n913 ); 
nand ( n1509 , n1496 , n1508 ); 
nand ( n1510 , n780 , n1509 ); 
nand ( n1511 , n1491 , n1510 ); 
and ( n1512 , n163 , n349 ); 
not ( n1513 , n348 ); 
or ( n1514 , n1512 , n1513 , n702 ); 
not ( n1515 , n347 ); 
or ( n1516 , n348 , n1515 , n16 ); 
nand ( n1517 , n1514 , n1516 ); 
not ( n1518 , n715 ); 
nand ( n1519 , n1518 , n708 ); 
not ( n1520 , n715 ); 
not ( n1521 , n733 ); 
nand ( n1522 , n345 , n1521 ); 
not ( n1523 , n1522 ); 
or ( n1524 , n1520 , n1523 ); 
nand ( n1525 , n1524 , n735 ); 
and ( n1526 , n1519 , n1525 ); 
nor ( n1527 , n1526 , n747 ); 
not ( n1528 , n256 ); 
not ( n1529 , n754 ); 
or ( n1530 , n1528 , n1529 ); 
nand ( n1531 , n257 , n758 ); 
nand ( n1532 , n1530 , n1531 ); 
nand ( n1533 , n258 , n763 ); 
nand ( n1534 , n260 , n766 ); 
nand ( n1535 , n259 , n771 ); 
nand ( n1536 , n1533 , n1534 , n1535 ); 
nor ( n1537 , n1532 , n1536 ); 
or ( n1538 , n1537 , n778 ); 
nand ( n1539 , n261 , n1163 ); 
nand ( n1540 , n262 , n1166 ); 
and ( n1541 , n1539 , n1540 ); 
nor ( n1542 , n1541 , n801 ); 
not ( n1543 , n1542 ); 
not ( n1544 , n263 ); 
not ( n1545 , n818 ); 
or ( n1546 , n1544 , n1545 ); 
nand ( n1547 , n266 , n841 ); 
nand ( n1548 , n1546 , n1547 ); 
not ( n1549 , n264 ); 
not ( n1550 , n834 ); 
or ( n1551 , n1549 , n1550 ); 
nand ( n1552 , n265 , n877 ); 
nand ( n1553 , n1551 , n1552 ); 
or ( n1554 , n1548 , n1553 ); 
nand ( n1555 , n1554 , n913 ); 
nand ( n1556 , n1543 , n1555 ); 
nand ( n1557 , n778 , n1556 ); 
nand ( n1558 , n1538 , n1557 ); 
and ( n1559 , n161 , n349 ); 
or ( n1560 , n1559 , n1513 , n652 ); 
not ( n1561 , n367 ); 
or ( n1562 , n1561 , n16 , n348 ); 
nand ( n1563 , n1560 , n1562 ); 
not ( n1564 , n801 ); 
and ( n1565 , n38 , n796 ); 
not ( n1566 , n14 ); 
not ( n1567 , n1052 ); 
or ( n1568 , n1566 , n1567 ); 
not ( n1569 , n790 ); 
nand ( n1570 , n37 , n1569 ); 
nand ( n1571 , n1568 , n1570 ); 
nor ( n1572 , n1565 , n1571 ); 
and ( n1573 , n1564 , n1572 ); 
not ( n1574 , n1564 ); 
not ( n1575 , n41 ); 
not ( n1576 , n834 ); 
or ( n1577 , n1575 , n1576 ); 
nand ( n1578 , n42 , n818 ); 
nand ( n1579 , n1577 , n1578 ); 
not ( n1580 , n40 ); 
not ( n1581 , n942 ); 
or ( n1582 , n1580 , n1581 ); 
nand ( n1583 , n39 , n824 ); 
nand ( n1584 , n1582 , n1583 ); 
nor ( n1585 , n1579 , n1584 ); 
and ( n1586 , n1574 , n1585 ); 
or ( n1587 , n1573 , n1586 ); 
and ( n1588 , n780 , n1587 ); 
not ( n1589 , n780 ); 
and ( n1590 , n34 , n771 ); 
and ( n1591 , n33 , n763 ); 
nor ( n1592 , n1590 , n1591 ); 
and ( n1593 , n31 , n754 ); 
and ( n1594 , n32 , n758 ); 
nor ( n1595 , n1593 , n1594 ); 
not ( n1596 , n1046 ); 
nand ( n1597 , n1596 , n35 , n1044 ); 
nand ( n1598 , n36 , n765 ); 
and ( n1599 , n1597 , n1598 ); 
nor ( n1600 , n1599 , 1'b0 ); 
and ( n1601 , n1592 , n1595 , n1600 ); 
and ( n1602 , n1589 , n1601 ); 
nor ( n1603 , n1588 , n1602 ); 
and ( n1604 , n201 , n1166 ); 
and ( n1605 , n72 , n1211 ); 
nor ( n1606 , n1604 , n1605 ); 
and ( n1607 , n1564 , n1606 ); 
not ( n1608 , n1564 ); 
not ( n1609 , n203 ); 
not ( n1610 , n834 ); 
or ( n1611 , n1609 , n1610 ); 
nand ( n1612 , n205 , n942 ); 
nand ( n1613 , n1611 , n1612 ); 
not ( n1614 , n202 ); 
not ( n1615 , n818 ); 
or ( n1616 , n1614 , n1615 ); 
nand ( n1617 , n204 , n824 ); 
nand ( n1618 , n1616 , n1617 ); 
nor ( n1619 , n1613 , n1618 ); 
and ( n1620 , n1608 , n1619 ); 
or ( n1621 , n1607 , n1620 ); 
and ( n1622 , n780 , n1621 ); 
not ( n1623 , n780 ); 
nand ( n1624 , n196 , n1047 ); 
nand ( n1625 , n198 , n763 ); 
nand ( n1626 , n197 , n852 ); 
nand ( n1627 , n1624 , n1625 , n1626 ); 
nand ( n1628 , n200 , n758 ); 
nand ( n1629 , n199 , n754 ); 
nand ( n1630 , n194 , n771 ); 
nand ( n1631 , n595 , n1234 ); 
nand ( n1632 , n1628 , n1629 , n1630 , n1631 ); 
nor ( n1633 , n1627 , n1632 ); 
and ( n1634 , n1623 , n1633 ); 
nor ( n1635 , n1622 , n1634 ); 
and ( n1636 , n239 , n1166 ); 
and ( n1637 , n14 , n1211 ); 
nor ( n1638 , n1636 , n1637 ); 
and ( n1639 , n1564 , n1638 ); 
not ( n1640 , n1564 ); 
not ( n1641 , n242 ); 
not ( n1642 , n818 ); 
or ( n1643 , n1641 , n1642 ); 
nand ( n1644 , n240 , n824 ); 
nand ( n1645 , n1643 , n1644 ); 
not ( n1646 , n243 ); 
not ( n1647 , n834 ); 
or ( n1648 , n1646 , n1647 ); 
nand ( n1649 , n241 , n841 ); 
nand ( n1650 , n1648 , n1649 ); 
nor ( n1651 , n1645 , n1650 ); 
and ( n1652 , n1640 , n1651 ); 
or ( n1653 , n1639 , n1652 ); 
and ( n1654 , n780 , n1653 ); 
not ( n1655 , n780 ); 
nand ( n1656 , n234 , n1047 ); 
nand ( n1657 , n238 , n763 ); 
nand ( n1658 , n237 , n852 ); 
nand ( n1659 , n1656 , n1657 , n1658 ); 
nand ( n1660 , n236 , n758 ); 
nand ( n1661 , n235 , n754 ); 
nand ( n1662 , n232 , n771 ); 
nand ( n1663 , n618 , n1234 ); 
nand ( n1664 , n1660 , n1661 , n1662 , n1663 ); 
nor ( n1665 , n1659 , n1664 ); 
and ( n1666 , n1655 , n1665 ); 
nor ( n1667 , n1654 , n1666 ); 
not ( n1668 , n801 ); 
and ( n1669 , n227 , n1166 ); 
and ( n1670 , n226 , n1211 ); 
nor ( n1671 , n1669 , n1670 ); 
and ( n1672 , n1668 , n1671 ); 
not ( n1673 , n1668 ); 
not ( n1674 , n229 ); 
not ( n1675 , n834 ); 
or ( n1676 , n1674 , n1675 ); 
nand ( n1677 , n228 , n818 ); 
nand ( n1678 , n1676 , n1677 ); 
not ( n1679 , n231 ); 
not ( n1680 , n942 ); 
or ( n1681 , n1679 , n1680 ); 
nand ( n1682 , n230 , n824 ); 
nand ( n1683 , n1681 , n1682 ); 
nor ( n1684 , n1678 , n1683 ); 
and ( n1685 , n1673 , n1684 ); 
or ( n1686 , n1672 , n1685 ); 
and ( n1687 , n780 , n1686 ); 
not ( n1688 , n780 ); 
nand ( n1689 , n221 , n1044 , n1047 ); 
nand ( n1690 , n223 , n763 ); 
nand ( n1691 , n222 , n852 ); 
nand ( n1692 , n1689 , n1690 , n1691 ); 
nand ( n1693 , n225 , n758 ); 
nand ( n1694 , n224 , n754 ); 
nand ( n1695 , n219 , n771 ); 
or ( n1696 , n16 , n220 ); 
nand ( n1697 , n1696 , n1234 ); 
nand ( n1698 , n1693 , n1694 , n1695 , n1697 ); 
nor ( n1699 , n1692 , n1698 ); 
and ( n1700 , n1688 , n1699 ); 
nor ( n1701 , n1687 , n1700 ); 
and ( n1702 , n214 , n1166 ); 
and ( n1703 , n213 , n1211 ); 
nor ( n1704 , n1702 , n1703 ); 
and ( n1705 , n1564 , n1704 ); 
not ( n1706 , n1564 ); 
not ( n1707 , n215 ); 
not ( n1708 , n834 ); 
or ( n1709 , n1707 , n1708 ); 
nand ( n1710 , n217 , n818 ); 
nand ( n1711 , n1709 , n1710 ); 
not ( n1712 , n216 ); 
not ( n1713 , n942 ); 
or ( n1714 , n1712 , n1713 ); 
nand ( n1715 , n218 , n824 ); 
nand ( n1716 , n1714 , n1715 ); 
nor ( n1717 , n1711 , n1716 ); 
and ( n1718 , n1706 , n1717 ); 
or ( n1719 , n1705 , n1718 ); 
and ( n1720 , n778 , n1719 ); 
not ( n1721 , n778 ); 
nand ( n1722 , n208 , n1047 ); 
nand ( n1723 , n210 , n763 ); 
nand ( n1724 , n209 , n852 ); 
nand ( n1725 , n1722 , n1723 , n1724 ); 
nand ( n1726 , n212 , n758 ); 
nand ( n1727 , n211 , n754 ); 
nand ( n1728 , n206 , n771 ); 
nand ( n1729 , n641 , n1234 ); 
nand ( n1730 , n1726 , n1727 , n1728 , n1729 ); 
nor ( n1731 , n1725 , n1730 ); 
and ( n1732 , n1721 , n1731 ); 
nor ( n1733 , n1720 , n1732 ); 
and ( n1734 , n295 , n1166 ); 
and ( n1735 , n48 , n1211 ); 
nor ( n1736 , n1734 , n1735 ); 
and ( n1737 , n1564 , n1736 ); 
not ( n1738 , n1564 ); 
not ( n1739 , n298 ); 
not ( n1740 , n834 ); 
or ( n1741 , n1739 , n1740 ); 
nand ( n1742 , n296 , n818 ); 
nand ( n1743 , n1741 , n1742 ); 
not ( n1744 , n297 ); 
not ( n1745 , n942 ); 
or ( n1746 , n1744 , n1745 ); 
nand ( n1747 , n299 , n824 ); 
nand ( n1748 , n1746 , n1747 ); 
nor ( n1749 , n1743 , n1748 ); 
and ( n1750 , n1738 , n1749 ); 
or ( n1751 , n1737 , n1750 ); 
and ( n1752 , n780 , n1751 ); 
not ( n1753 , n780 ); 
nand ( n1754 , n291 , n1047 ); 
nand ( n1755 , n294 , n763 ); 
nand ( n1756 , n293 , n852 ); 
nand ( n1757 , n1754 , n1755 , n1756 ); 
nand ( n1758 , n292 , n758 ); 
nand ( n1759 , n156 , n754 ); 
nand ( n1760 , n289 , n771 ); 
nand ( n1761 , n554 , n1234 ); 
nand ( n1762 , n1758 , n1759 , n1760 , n1761 ); 
nor ( n1763 , n1757 , n1762 ); 
and ( n1764 , n1753 , n1763 ); 
nor ( n1765 , n1752 , n1764 ); 
not ( n1766 , n345 ); 
not ( n1767 , n717 ); 
and ( n1768 , n1766 , n1767 ); 
not ( n1769 , n345 ); 
not ( n1770 , n732 ); 
or ( n1771 , n1769 , n1770 ); 
nand ( n1772 , n1771 , n717 ); 
and ( n1773 , n733 , n1772 ); 
nor ( n1774 , n1768 , n1773 ); 
nor ( n1775 , n747 , n1774 ); 
nand ( n1776 , n708 , n720 ); 
not ( n1777 , n732 ); 
nor ( n1778 , n725 , n730 ); 
nand ( n1779 , n1777 , t_0 , n345 ); 
and ( n1780 , n1776 , n1779 ); 
nor ( n1781 , n1780 , n747 ); 
not ( n1782 , n1597 ); 
not ( n1783 , n338 ); 
nor ( n1784 , n341 , n342 ); 
not ( n1785 , n339 ); 
nor ( n1786 , n1785 , n340 ); 
not ( n1787 , n153 ); 
nor ( n1788 , n1787 , n16 ); 
nand ( n1789 , n1783 , n1784 , n1786 , n1788 ); 
not ( n1790 , n1789 ); 
or ( n1791 , n278 , n1790 ); 
nor ( n1792 , n16 , n343 ); 
not ( n1793 , n160 ); 
nand ( n1794 , n1793 , n1790 ); 
nand ( n1795 , n1791 , n1792 , n1794 ); 
not ( n1796 , n1792 ); 
nand ( n1797 , n289 , n1796 ); 
nand ( n1798 , n317 , n1796 ); 
nand ( n1799 , n1795 , n1797 , n1798 ); 
nand ( n1800 , n708 , n723 ); 
or ( n1801 , n722 , n1778 ); 
nand ( n1802 , n722 , n1778 ); 
nand ( n1803 , n1801 , n1802 , n345 ); 
and ( n1804 , n1800 , n1803 ); 
nor ( n1805 , n1804 , n747 ); 
and ( n1806 , n337 , n1790 ); 
and ( n1807 , n247 , n1789 ); 
nor ( n1808 , n1806 , n1807 ); 
or ( n1809 , n1796 , n1808 ); 
nand ( n1810 , n1809 , n1798 ); 
and ( n1811 , n336 , n1790 ); 
and ( n1812 , n312 , n1789 ); 
nor ( n1813 , n1811 , n1812 ); 
or ( n1814 , n1796 , n1813 ); 
nand ( n1815 , n1814 , n1797 ); 
not ( n1816 , n345 ); 
not ( n1817 , n729 ); 
not ( n1818 , n1817 ); 
and ( n1819 , n1816 , n1818 ); 
not ( n1820 , n727 ); 
and ( n1821 , n1820 , n1817 ); 
nand ( n1822 , n345 , n730 ); 
nor ( n1823 , n1821 , n1822 ); 
nor ( n1824 , n1819 , n1823 ); 
nor ( n1825 , n747 , n1824 ); 
not ( n1826 , n1778 ); 
or ( n1827 , n708 , n730 ); 
nand ( n1828 , n1827 , n725 ); 
and ( n1829 , n1826 , n1828 ); 
not ( n1830 , n725 ); 
and ( n1831 , n708 , n1830 ); 
nor ( n1832 , n1829 , n1831 ); 
nor ( n1833 , n747 , n1832 ); 
nor ( n1834 , n154 , n155 ); 
not ( n1835 , n151 ); 
nor ( n1836 , n1835 , n152 ); 
nand ( n1837 , n1834 , n1836 , n150 , n1788 ); 
nand ( n1838 , n249 , n1837 ); 
not ( n1839 , n1837 ); 
nand ( n1840 , n337 , n1839 ); 
and ( n1841 , n1838 , n1840 ); 
or ( n1842 , n16 , n158 ); 
nor ( n1843 , n1841 , n1842 ); 
nand ( n1844 , n314 , n1837 ); 
nand ( n1845 , n336 , n1839 ); 
and ( n1846 , n1844 , n1845 ); 
nor ( n1847 , n1846 , n1842 ); 
nand ( n1848 , n156 , n1837 ); 
nand ( n1849 , n157 , n1839 ); 
and ( n1850 , n1848 , n1849 ); 
nor ( n1851 , n1850 , n1842 ); 
nand ( n1852 , n159 , n1837 ); 
nand ( n1853 , n160 , n1839 ); 
and ( n1854 , n1852 , n1853 ); 
nor ( n1855 , n1854 , n1842 ); 
and ( n1856 , n1790 , n157 ); 
not ( n1857 , n1790 ); 
and ( n1858 , n1857 , n293 ); 
nor ( n1859 , n1856 , n1858 ); 
nor ( n1860 , n1796 , n1859 ); 
not ( n1861 , n1018 ); 
not ( n1862 , n1021 ); 
not ( n1863 , n1598 ); 
and ( n1864 , n345 , n1820 , n746 ); 
and ( n1865 , n374 , n1044 ); 
nor ( n1866 , n1865 , n373 ); 
nor ( n1867 , n747 , n1866 ); 
not ( n1868 , n379 ); 
not ( n1869 , n16 ); 
nand ( n1870 , n1869 , n378 ); 
nand ( n1871 , n1868 , n1870 ); 
nor ( n1872 , n376 , n377 ); 
nor ( n1873 , n16 , n1872 ); 
and ( n1874 , n371 , n351 ); 
not ( n1875 , n371 ); 
and ( n1876 , n1875 , n389 ); 
or ( n1877 , n1874 , n1876 ); 
and ( n1878 , n371 , n386 ); 
not ( n1879 , n371 ); 
and ( n1880 , n1879 , n385 ); 
or ( n1881 , n1878 , n1880 ); 
and ( n1882 , n371 , n393 ); 
not ( n1883 , n371 ); 
and ( n1884 , n1883 , n392 ); 
or ( n1885 , n1882 , n1884 ); 
and ( n1886 , n371 , n400 ); 
not ( n1887 , n371 ); 
and ( n1888 , n1887 , n399 ); 
or ( n1889 , n1886 , n1888 ); 
and ( n1890 , n371 , n354 ); 
not ( n1891 , n371 ); 
and ( n1892 , n1891 , n390 ); 
or ( n1893 , n1890 , n1892 ); 
and ( n1894 , n371 , n4 ); 
not ( n1895 , n371 ); 
and ( n1896 , n1895 , n394 ); 
or ( n1897 , n1894 , n1896 ); 
and ( n1898 , n371 , n388 ); 
not ( n1899 , n371 ); 
and ( n1900 , n1899 , n387 ); 
or ( n1901 , n1898 , n1900 ); 
and ( n1902 , n371 , n407 ); 
not ( n1903 , n371 ); 
and ( n1904 , n1903 , n406 ); 
or ( n1905 , n1902 , n1904 ); 
and ( n1906 , n371 , n398 ); 
not ( n1907 , n371 ); 
and ( n1908 , n1907 , n397 ); 
or ( n1909 , n1906 , n1908 ); 
and ( n1910 , n371 , n405 ); 
not ( n1911 , n371 ); 
and ( n1912 , n1911 , n404 ); 
or ( n1913 , n1910 , n1912 ); 
and ( n1914 , n371 , n2 ); 
not ( n1915 , n371 ); 
and ( n1916 , n1915 , n403 ); 
or ( n1917 , n1914 , n1916 ); 
and ( n1918 , n371 , n3 ); 
not ( n1919 , n371 ); 
and ( n1920 , n1919 , n391 ); 
or ( n1921 , n1918 , n1920 ); 
and ( n1922 , n371 , n396 ); 
not ( n1923 , n371 ); 
and ( n1924 , n1923 , n395 ); 
or ( n1925 , n1922 , n1924 ); 
and ( n1926 , n371 , n6 ); 
not ( n1927 , n371 ); 
and ( n1928 , n1927 , n408 ); 
or ( n1929 , n1926 , n1928 ); 
and ( n1930 , n371 , n5 ); 
not ( n1931 , n371 ); 
and ( n1932 , n1931 , n411 ); 
or ( n1933 , n1930 , n1932 ); 
and ( n1934 , n371 , n410 ); 
not ( n1935 , n371 ); 
and ( n1936 , n1935 , n409 ); 
or ( n1937 , n1934 , n1936 ); 
and ( n1938 , n371 , n402 ); 
not ( n1939 , n371 ); 
and ( n1940 , n1939 , n401 ); 
or ( n1941 , n1938 , n1940 ); 
or ( n1942 , n16 , n382 ); 
not ( n1943 , n375 ); 
nor ( n1944 , n1943 , n16 ); 
or ( n1945 , n16 , n383 ); 
or ( n1946 , n16 , n380 ); 
or ( n1947 , n16 , n381 ); 
or ( n1948 , n16 , n384 ); 
patch p0 (.t_0(t_0), .g1(n1778), .g2(n1805), .g3(n720));
endmodule 

