module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 ; 
output g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 ; 
wire t_0 , t_1 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( n158 , g157 ); 
buf ( n159 , g158 ); 
buf ( n160 , g159 ); 
buf ( n161 , g160 ); 
buf ( n162 , g161 ); 
buf ( n163 , g162 ); 
buf ( n164 , g163 ); 
buf ( n165 , g164 ); 
buf ( n166 , g165 ); 
buf ( n167 , g166 ); 
buf ( n168 , g167 ); 
buf ( n169 , g168 ); 
buf ( n170 , g169 ); 
buf ( n171 , g170 ); 
buf ( n172 , g171 ); 
buf ( n173 , g172 ); 
buf ( n174 , g173 ); 
buf ( n175 , g174 ); 
buf ( n176 , g175 ); 
buf ( n177 , g176 ); 
buf ( n178 , g177 ); 
buf ( n179 , g178 ); 
buf ( n180 , g179 ); 
buf ( n181 , g180 ); 
buf ( n182 , g181 ); 
buf ( n183 , g182 ); 
buf ( n184 , g183 ); 
buf ( n185 , g184 ); 
buf ( n186 , g185 ); 
buf ( n187 , g186 ); 
buf ( n188 , g187 ); 
buf ( n189 , g188 ); 
buf ( n190 , g189 ); 
buf ( n191 , g190 ); 
buf ( n192 , g191 ); 
buf ( n193 , g192 ); 
buf ( n194 , g193 ); 
buf ( n195 , g194 ); 
buf ( n196 , g195 ); 
buf ( n197 , g196 ); 
buf ( n198 , g197 ); 
buf ( n199 , g198 ); 
buf ( n200 , g199 ); 
buf ( n201 , g200 ); 
buf ( n202 , g201 ); 
buf ( n203 , g202 ); 
buf ( n204 , g203 ); 
buf ( n205 , g204 ); 
buf ( n206 , g205 ); 
buf ( n207 , g206 ); 
buf ( n208 , g207 ); 
buf ( n209 , g208 ); 
buf ( n210 , g209 ); 
buf ( n211 , g210 ); 
buf ( n212 , g211 ); 
buf ( n213 , g212 ); 
buf ( n214 , g213 ); 
buf ( n215 , g214 ); 
buf ( n216 , g215 ); 
buf ( n217 , g216 ); 
buf ( n218 , g217 ); 
buf ( n219 , g218 ); 
buf ( n220 , g219 ); 
buf ( n221 , g220 ); 
buf ( n222 , g221 ); 
buf ( n223 , g222 ); 
buf ( n224 , g223 ); 
buf ( n225 , g224 ); 
buf ( n226 , g225 ); 
buf ( n227 , g226 ); 
buf ( n228 , g227 ); 
buf ( n229 , g228 ); 
buf ( n230 , g229 ); 
buf ( n231 , g230 ); 
buf ( n232 , g231 ); 
buf ( n233 , g232 ); 
buf ( n234 , g233 ); 
buf ( n235 , g234 ); 
buf ( n236 , g235 ); 
buf ( n237 , g236 ); 
buf ( n238 , g237 ); 
buf ( n239 , g238 ); 
buf ( n240 , g239 ); 
buf ( n241 , g240 ); 
buf ( n242 , g241 ); 
buf ( n243 , g242 ); 
buf ( n244 , g243 ); 
buf ( n245 , g244 ); 
buf ( n246 , g245 ); 
buf ( n247 , g246 ); 
buf ( n248 , g247 ); 
buf ( n249 , g248 ); 
buf ( n250 , g249 ); 
buf ( n251 , g250 ); 
buf ( n252 , g251 ); 
buf ( n253 , g252 ); 
buf ( n254 , g253 ); 
buf ( n255 , g254 ); 
buf ( n256 , g255 ); 
buf ( n257 , g256 ); 
buf ( n258 , g257 ); 
buf ( n259 , g258 ); 
buf ( n260 , g259 ); 
buf ( n261 , g260 ); 
buf ( n262 , g261 ); 
buf ( n263 , g262 ); 
buf ( n264 , g263 ); 
buf ( n265 , g264 ); 
buf ( n266 , g265 ); 
buf ( n267 , g266 ); 
buf ( n268 , g267 ); 
buf ( n269 , g268 ); 
buf ( n270 , g269 ); 
buf ( n271 , g270 ); 
buf ( n272 , g271 ); 
buf ( n273 , g272 ); 
buf ( n274 , g273 ); 
buf ( n275 , g274 ); 
buf ( n276 , g275 ); 
buf ( n277 , g276 ); 
buf ( n278 , g277 ); 
buf ( n279 , g278 ); 
buf ( n280 , g279 ); 
buf ( n281 , g280 ); 
buf ( n282 , g281 ); 
buf ( n283 , g282 ); 
buf ( n284 , g283 ); 
buf ( n285 , g284 ); 
buf ( n286 , g285 ); 
buf ( n287 , g286 ); 
buf ( n288 , g287 ); 
buf ( n289 , g288 ); 
buf ( n290 , g289 ); 
buf ( n291 , g290 ); 
buf ( n292 , g291 ); 
buf ( n293 , g292 ); 
buf ( n294 , g293 ); 
buf ( n295 , g294 ); 
buf ( n296 , g295 ); 
buf ( n297 , g296 ); 
buf ( n298 , g297 ); 
buf ( n299 , g298 ); 
buf ( n300 , g299 ); 
buf ( n301 , g300 ); 
buf ( n302 , g301 ); 
buf ( n303 , g302 ); 
buf ( n304 , g303 ); 
buf ( n305 , g304 ); 
buf ( n306 , g305 ); 
buf ( n307 , g306 ); 
buf ( n308 , g307 ); 
buf ( n309 , g308 ); 
buf ( n310 , g309 ); 
buf ( n311 , g310 ); 
buf ( n312 , g311 ); 
buf ( n313 , g312 ); 
buf ( n314 , g313 ); 
buf ( n315 , g314 ); 
buf ( n316 , g315 ); 
buf ( n317 , g316 ); 
buf ( n318 , g317 ); 
buf ( n319 , g318 ); 
buf ( n320 , g319 ); 
buf ( n321 , g320 ); 
buf ( n322 , g321 ); 
buf ( n323 , g322 ); 
buf ( n324 , g323 ); 
buf ( n325 , g324 ); 
buf ( n326 , g325 ); 
buf ( n327 , g326 ); 
buf ( n328 , g327 ); 
buf ( n329 , g328 ); 
buf ( n330 , g329 ); 
buf ( n331 , g330 ); 
buf ( n332 , g331 ); 
buf ( n333 , g332 ); 
buf ( n334 , g333 ); 
buf ( n335 , g334 ); 
buf ( n336 , g335 ); 
buf ( n337 , g336 ); 
buf ( n338 , g337 ); 
buf ( n339 , g338 ); 
buf ( n340 , g339 ); 
buf ( n341 , g340 ); 
buf ( n342 , g341 ); 
buf ( n343 , g342 ); 
buf ( n344 , g343 ); 
buf ( n345 , g344 ); 
buf ( n346 , g345 ); 
buf ( n347 , g346 ); 
buf ( n348 , g347 ); 
buf ( n349 , g348 ); 
buf ( n350 , g349 ); 
buf ( n351 , g350 ); 
buf ( n352 , g351 ); 
buf ( n353 , g352 ); 
buf ( n354 , g353 ); 
buf ( n355 , g354 ); 
buf ( n356 , g355 ); 
buf ( n357 , g356 ); 
buf ( n358 , g357 ); 
buf ( n359 , g358 ); 
buf ( n360 , g359 ); 
buf ( n361 , g360 ); 
buf ( n362 , g361 ); 
buf ( n363 , g362 ); 
buf ( n364 , g363 ); 
buf ( n365 , g364 ); 
buf ( n366 , g365 ); 
buf ( n367 , g366 ); 
buf ( n368 , g367 ); 
buf ( n369 , g368 ); 
buf ( n370 , g369 ); 
buf ( n371 , g370 ); 
buf ( n372 , g371 ); 
buf ( n373 , g372 ); 
buf ( n374 , g373 ); 
buf ( n375 , g374 ); 
buf ( n376 , g375 ); 
buf ( n377 , g376 ); 
buf ( n378 , g377 ); 
buf ( n379 , g378 ); 
buf ( n380 , g379 ); 
buf ( n381 , g380 ); 
buf ( n382 , g381 ); 
buf ( n383 , g382 ); 
buf ( n384 , g383 ); 
buf ( n385 , g384 ); 
buf ( n386 , g385 ); 
buf ( n387 , g386 ); 
buf ( n388 , g387 ); 
buf ( n389 , g388 ); 
buf ( n390 , g389 ); 
buf ( n391 , g390 ); 
buf ( n392 , g391 ); 
buf ( n393 , g392 ); 
buf ( n394 , g393 ); 
buf ( n395 , g394 ); 
buf ( n396 , g395 ); 
buf ( n397 , g396 ); 
buf ( n398 , g397 ); 
buf ( n399 , g398 ); 
buf ( n400 , g399 ); 
buf ( n401 , g400 ); 
buf ( n402 , g401 ); 
buf ( n403 , g402 ); 
buf ( n404 , g403 ); 
buf ( n405 , g404 ); 
buf ( n406 , g405 ); 
buf ( n407 , g406 ); 
buf ( n408 , g407 ); 
buf ( n409 , g408 ); 
buf ( n410 , g409 ); 
buf ( n411 , g410 ); 
buf ( n412 , g411 ); 
buf ( n413 , g412 ); 
buf ( n414 , g413 ); 
buf ( n415 , g414 ); 
buf ( n416 , g415 ); 
buf ( n417 , g416 ); 
buf ( g417 , n418 ); 
buf ( g418 , n419 ); 
buf ( g419 , n420 ); 
buf ( g420 , n421 ); 
buf ( g421 , n422 ); 
buf ( g422 , n423 ); 
buf ( g423 , n424 ); 
buf ( g424 , n425 ); 
buf ( g425 , n426 ); 
buf ( g426 , n427 ); 
buf ( g427 , n428 ); 
buf ( g428 , n429 ); 
buf ( g429 , n430 ); 
buf ( g430 , n431 ); 
buf ( g431 , n432 ); 
buf ( g432 , n433 ); 
buf ( g433 , n434 ); 
buf ( g434 , n435 ); 
buf ( g435 , n436 ); 
buf ( g436 , n437 ); 
buf ( g437 , n438 ); 
buf ( g438 , n439 ); 
buf ( g439 , n440 ); 
buf ( g440 , n441 ); 
buf ( g441 , n442 ); 
buf ( g442 , n443 ); 
buf ( g443 , n444 ); 
buf ( g444 , n445 ); 
buf ( g445 , n446 ); 
buf ( g446 , n447 ); 
buf ( g447 , n448 ); 
buf ( g448 , n449 ); 
buf ( g449 , n450 ); 
buf ( g450 , n451 ); 
buf ( g451 , n452 ); 
buf ( g452 , n453 ); 
buf ( g453 , n454 ); 
buf ( g454 , n455 ); 
buf ( g455 , n456 ); 
buf ( g456 , n457 ); 
buf ( g457 , n458 ); 
buf ( g458 , n459 ); 
buf ( g459 , n460 ); 
buf ( g460 , n461 ); 
buf ( g461 , n462 ); 
buf ( g462 , n463 ); 
buf ( g463 , n464 ); 
buf ( g464 , n465 ); 
buf ( g465 , n466 ); 
buf ( g466 , n467 ); 
buf ( g467 , n468 ); 
buf ( g468 , n469 ); 
buf ( g469 , n470 ); 
buf ( g470 , n471 ); 
buf ( g471 , n472 ); 
buf ( g472 , n473 ); 
buf ( g473 , n474 ); 
buf ( g474 , n475 ); 
buf ( g475 , n476 ); 
buf ( g476 , n477 ); 
buf ( g477 , n478 ); 
buf ( g478 , n479 ); 
buf ( g479 , n480 ); 
buf ( g480 , n481 ); 
buf ( g481 , n482 ); 
buf ( g482 , n483 ); 
buf ( g483 , n484 ); 
buf ( g484 , n485 ); 
buf ( g485 , n486 ); 
buf ( g486 , n487 ); 
buf ( g487 , n488 ); 
buf ( g488 , n489 ); 
buf ( g489 , n490 ); 
buf ( g490 , n491 ); 
buf ( g491 , n492 ); 
buf ( g492 , n493 ); 
buf ( g493 , n494 ); 
buf ( g494 , n495 ); 
buf ( g495 , n496 ); 
buf ( g496 , n497 ); 
buf ( g497 , n498 ); 
buf ( g498 , n499 ); 
buf ( g499 , n500 ); 
buf ( g500 , n501 ); 
buf ( g501 , n502 ); 
buf ( g502 , n503 ); 
buf ( g503 , n504 ); 
buf ( g504 , n505 ); 
buf ( g505 , n506 ); 
buf ( g506 , n507 ); 
buf ( g507 , n508 ); 
buf ( g508 , n509 ); 
buf ( g509 , n510 ); 
buf ( g510 , n511 ); 
buf ( g511 , n512 ); 
buf ( g512 , n513 ); 
buf ( g513 , n514 ); 
buf ( g514 , n515 ); 
buf ( g515 , n516 ); 
buf ( g516 , n517 ); 
buf ( g517 , n518 ); 
buf ( g518 , n519 ); 
buf ( g519 , n520 ); 
buf ( g520 , n521 ); 
buf ( g521 , n522 ); 
buf ( g522 , n523 ); 
buf ( g523 , n524 ); 
buf ( g524 , n525 ); 
buf ( g525 , n526 ); 
buf ( g526 , n527 ); 
buf ( g527 , n528 ); 
buf ( g528 , n529 ); 
buf ( g529 , n530 ); 
buf ( g530 , n531 ); 
buf ( g531 , n532 ); 
buf ( g532 , n533 ); 
buf ( g533 , n534 ); 
buf ( g534 , n535 ); 
buf ( g535 , n536 ); 
buf ( g536 , n537 ); 
buf ( g537 , n538 ); 
buf ( g538 , n539 ); 
buf ( g539 , n540 ); 
buf ( g540 , n541 ); 
buf ( g541 , n542 ); 
buf ( g542 , n543 ); 
buf ( g543 , n544 ); 
buf ( g544 , n545 ); 
buf ( g545 , n546 ); 
buf ( g546 , n547 ); 
buf ( g547 , n548 ); 
buf ( g548 , n549 ); 
buf ( g549 , n550 ); 
buf ( g550 , n551 ); 
buf ( g551 , n552 ); 
buf ( g552 , n553 ); 
buf ( g553 , n554 ); 
buf ( g554 , n555 ); 
buf ( g555 , n556 ); 
buf ( g556 , n557 ); 
buf ( g557 , n558 ); 
buf ( g558 , n559 ); 
buf ( g559 , n560 ); 
buf ( g560 , n561 ); 
buf ( g561 , n562 ); 
buf ( g562 , n563 ); 
buf ( g563 , n564 ); 
buf ( g564 , n565 ); 
buf ( g565 , n566 ); 
buf ( g566 , n567 ); 
buf ( g567 , n568 ); 
buf ( g568 , n569 ); 
buf ( g569 , n570 ); 
buf ( g570 , n571 ); 
buf ( g571 , n572 ); 
buf ( g572 , n573 ); 
buf ( g573 , n574 ); 
buf ( g574 , n575 ); 
buf ( g575 , n576 ); 
buf ( g576 , n577 ); 
buf ( g577 , n578 ); 
buf ( g578 , n579 ); 
buf ( g579 , n580 ); 
buf ( g580 , n581 ); 
buf ( g581 , n582 ); 
buf ( g582 , n583 ); 
buf ( g583 , n584 ); 
buf ( g584 , n585 ); 
buf ( g585 , n586 ); 
buf ( g586 , n587 ); 
buf ( g587 , n588 ); 
buf ( g588 , n589 ); 
buf ( g589 , n590 ); 
buf ( g590 , n591 ); 
buf ( g591 , n592 ); 
buf ( g592 , n593 ); 
buf ( g593 , n594 ); 
buf ( g594 , n595 ); 
buf ( g595 , n596 ); 
buf ( g596 , n597 ); 
buf ( g597 , n598 ); 
buf ( g598 , n599 ); 
buf ( g599 , n600 ); 
buf ( g600 , n601 ); 
buf ( g601 , n602 ); 
buf ( g602 , n603 ); 
buf ( g603 , n604 ); 
buf ( g604 , n605 ); 
buf ( g605 , n606 ); 
buf ( g606 , n607 ); 
buf ( g607 , n608 ); 
buf ( g608 , n609 ); 
buf ( g609 , n610 ); 
buf ( g610 , n611 ); 
buf ( g611 , n612 ); 
buf ( g612 , n613 ); 
buf ( g613 , n614 ); 
buf ( g614 , n615 ); 
buf ( g615 , n616 ); 
buf ( g616 , n617 ); 
buf ( g617 , n618 ); 
buf ( g618 , n619 ); 
buf ( g619 , n620 ); 
buf ( g620 , n621 ); 
buf ( g621 , n622 ); 
buf ( g622 , n623 ); 
buf ( g623 , n624 ); 
buf ( g624 , n625 ); 
buf ( g625 , n626 ); 
buf ( g626 , n627 ); 
buf ( g627 , n628 ); 
buf ( g628 , n629 ); 
buf ( g629 , n630 ); 
buf ( g630 , n631 ); 
buf ( n418 , 1'b0 ); 
buf ( n419 , n2138 ); 
buf ( n420 , 1'b0 ); 
buf ( n421 , n2134 ); 
buf ( n422 , 1'b0 ); 
buf ( n423 , n2131 ); 
buf ( n424 , 1'b0 ); 
buf ( n425 , 1'b0 ); 
buf ( n426 , n2142 ); 
buf ( n427 , 1'b0 ); 
buf ( n428 , n2149 ); 
buf ( n429 , n2112 ); 
buf ( n430 , 1'b0 ); 
buf ( n431 , n2145 ); 
buf ( n432 , n1947 ); 
buf ( n433 , n2210 ); 
buf ( n434 , n2151 ); 
buf ( n435 , n2150 ); 
buf ( n436 , n1991 ); 
buf ( n437 , n1930 ); 
buf ( n438 , n2154 ); 
buf ( n439 , n2155 ); 
buf ( n440 , n2156 ); 
buf ( n441 , n1991 ); 
buf ( n442 , n2129 ); 
buf ( n443 , n2158 ); 
buf ( n444 , n2160 ); 
buf ( n445 , n1985 ); 
buf ( n446 , n2161 ); 
buf ( n447 , n2113 ); 
buf ( n448 , n2162 ); 
buf ( n449 , n2164 ); 
buf ( n450 , n2166 ); 
buf ( n451 , n2147 ); 
buf ( n452 , n2167 ); 
buf ( n453 , 1'b0 ); 
buf ( n454 , n2110 ); 
buf ( n455 , n2211 ); 
buf ( n456 , n2065 ); 
buf ( n457 , n2169 ); 
buf ( n458 , n2213 ); 
buf ( n459 , n2170 ); 
buf ( n460 , n2035 ); 
buf ( n461 , n2195 ); 
buf ( n462 , n2171 ); 
buf ( n463 , n2209 ); 
buf ( n464 , n2173 ); 
buf ( n465 , n2175 ); 
buf ( n466 , n2177 ); 
buf ( n467 , n2140 ); 
buf ( n468 , n2068 ); 
buf ( n469 , n2181 ); 
buf ( n470 , n1962 ); 
buf ( n471 , n2179 ); 
buf ( n472 , n2144 ); 
buf ( n473 , n2094 ); 
buf ( n474 , n2182 ); 
buf ( n475 , 1'b0 ); 
buf ( n476 , n2095 ); 
buf ( n477 , n2136 ); 
buf ( n478 , n2098 ); 
buf ( n479 , n2183 ); 
buf ( n480 , 1'b0 ); 
buf ( n481 , n2084 ); 
buf ( n482 , n2133 ); 
buf ( n483 , n2099 ); 
buf ( n484 , n2184 ); 
buf ( n485 , 1'b0 ); 
buf ( n486 , n2128 ); 
buf ( n487 , n2100 ); 
buf ( n488 , n2148 ); 
buf ( n489 , 1'b0 ); 
buf ( n490 , n2186 ); 
buf ( n491 , n2214 ); 
buf ( n492 , n2188 ); 
buf ( n493 , n2194 ); 
buf ( n494 , n2190 ); 
buf ( n495 , 1'b0 ); 
buf ( n496 , n2191 ); 
buf ( n497 , n2193 ); 
buf ( n498 , 1'b0 ); 
buf ( n499 , n2146 ); 
buf ( n500 , 1'b0 ); 
buf ( n501 , 1'b0 ); 
buf ( n502 , n1 ); 
buf ( n503 , n2236 ); 
buf ( n504 , 1'b0 ); 
buf ( n505 , 1'b0 ); 
buf ( n506 , n1 ); 
buf ( n507 , n1868 ); 
buf ( n508 , 1'b0 ); 
buf ( n509 , 1'b0 ); 
buf ( n510 , n1 ); 
buf ( n511 , n1680 ); 
buf ( n512 , 1'b0 ); 
buf ( n513 , 1'b0 ); 
buf ( n514 , n1 ); 
buf ( n515 , n1172 ); 
buf ( n516 , 1'b0 ); 
buf ( n517 , 1'b0 ); 
buf ( n518 , n1 ); 
buf ( n519 , n2034 ); 
buf ( n520 , 1'b0 ); 
buf ( n521 , 1'b0 ); 
buf ( n522 , n1 ); 
buf ( n523 , n1993 ); 
buf ( n524 , 1'b0 ); 
buf ( n525 , 1'b0 ); 
buf ( n526 , n1 ); 
buf ( n527 , n2108 ); 
buf ( n528 , 1'b0 ); 
buf ( n529 , 1'b0 ); 
buf ( n530 , n1 ); 
buf ( n531 , n1470 ); 
buf ( n532 , 1'b0 ); 
buf ( n533 , 1'b0 ); 
buf ( n534 , n1 ); 
buf ( n535 , n2025 ); 
buf ( n536 , 1'b0 ); 
buf ( n537 , 1'b0 ); 
buf ( n538 , n1 ); 
buf ( n539 , n1834 ); 
buf ( n540 , 1'b0 ); 
buf ( n541 , 1'b0 ); 
buf ( n542 , n1 ); 
buf ( n543 , n2234 ); 
buf ( n544 , 1'b0 ); 
buf ( n545 , 1'b0 ); 
buf ( n546 , n1 ); 
buf ( n547 , n1914 ); 
buf ( n548 , 1'b0 ); 
buf ( n549 , 1'b0 ); 
buf ( n550 , n1 ); 
buf ( n551 , n1734 ); 
buf ( n552 , 1'b0 ); 
buf ( n553 , 1'b0 ); 
buf ( n554 , n1 ); 
buf ( n555 , n2126 ); 
buf ( n556 , 1'b0 ); 
buf ( n557 , 1'b0 ); 
buf ( n558 , n1 ); 
buf ( n559 , n1998 ); 
buf ( n560 , 1'b0 ); 
buf ( n561 , 1'b0 ); 
buf ( n562 , n1 ); 
buf ( n563 , n1640 ); 
buf ( n564 , 1'b0 ); 
buf ( n565 , 1'b0 ); 
buf ( n566 , n1 ); 
buf ( n567 , n1955 ); 
buf ( n568 , 1'b0 ); 
buf ( n569 , 1'b0 ); 
buf ( n570 , n1 ); 
buf ( n571 , n2004 ); 
buf ( n572 , 1'b0 ); 
buf ( n573 , 1'b0 ); 
buf ( n574 , n1 ); 
buf ( n575 , n2092 ); 
buf ( n576 , 1'b0 ); 
buf ( n577 , 1'b0 ); 
buf ( n578 , n1 ); 
buf ( n579 , n2053 ); 
buf ( n580 , 1'b0 ); 
buf ( n581 , 1'b0 ); 
buf ( n582 , n1 ); 
buf ( n583 , n1572 ); 
buf ( n584 , 1'b0 ); 
buf ( n585 , 1'b0 ); 
buf ( n586 , n1 ); 
buf ( n587 , n1966 ); 
buf ( n588 , 1'b0 ); 
buf ( n589 , 1'b0 ); 
buf ( n590 , n1 ); 
buf ( n591 , n1936 ); 
buf ( n592 , 1'b0 ); 
buf ( n593 , 1'b0 ); 
buf ( n594 , n1 ); 
buf ( n595 , n2218 ); 
buf ( n596 , 1'b0 ); 
buf ( n597 , 1'b0 ); 
buf ( n598 , n1 ); 
buf ( n599 , n2228 ); 
buf ( n600 , 1'b0 ); 
buf ( n601 , 1'b0 ); 
buf ( n602 , n1 ); 
buf ( n603 , n2202 ); 
buf ( n604 , 1'b0 ); 
buf ( n605 , 1'b0 ); 
buf ( n606 , n1 ); 
buf ( n607 , n2208 ); 
buf ( n608 , 1'b0 ); 
buf ( n609 , 1'b0 ); 
buf ( n610 , n1 ); 
buf ( n611 , n2014 ); 
buf ( n612 , 1'b0 ); 
buf ( n613 , 1'b0 ); 
buf ( n614 , n1 ); 
buf ( n615 , n1988 ); 
buf ( n616 , 1'b0 ); 
buf ( n617 , 1'b0 ); 
buf ( n618 , n1 ); 
buf ( n619 , n2017 ); 
buf ( n620 , 1'b0 ); 
buf ( n621 , 1'b0 ); 
buf ( n622 , n1 ); 
buf ( n623 , n2067 ); 
buf ( n624 , 1'b0 ); 
buf ( n625 , 1'b0 ); 
buf ( n626 , n1 ); 
buf ( n627 , n1918 ); 
buf ( n628 , 1'b0 ); 
buf ( n629 , 1'b0 ); 
buf ( n630 , n1 ); 
buf ( n631 , n2223 ); 
and ( n714 , n388 , n401 ); 
nor ( n715 , n390 , n394 ); 
not ( n716 , n715 ); 
buf ( n717 , n716 ); 
not ( n718 , n344 ); 
nor ( n719 , n717 , n718 ); 
not ( n720 , n719 ); 
not ( n721 , n373 ); 
nand ( n722 , n721 , n359 ); 
nand ( n723 , n722 , n391 ); 
not ( n724 , n359 ); 
nor ( n725 , n724 , n373 ); 
nand ( n726 , n725 , n389 ); 
not ( n727 , n395 ); 
and ( n728 , n723 , n726 , n727 ); 
not ( n729 , n393 ); 
nand ( n730 , n729 , n359 ); 
and ( n731 , n728 , n730 ); 
not ( n732 , n731 ); 
not ( n733 , n732 ); 
or ( n734 , n720 , n733 ); 
nor ( n735 , n389 , n391 ); 
not ( n736 , n735 ); 
nand ( n737 , n717 , n736 , n398 ); 
nand ( n738 , n734 , n737 ); 
and ( n739 , n714 , n738 ); 
and ( n740 , n311 , n409 ); 
not ( n741 , n311 ); 
not ( n742 , n409 ); 
and ( n743 , n741 , n742 ); 
nor ( n744 , n740 , n743 ); 
not ( n745 , n744 ); 
and ( n746 , n413 , n24 ); 
not ( n747 , n413 ); 
and ( n748 , n747 , n64 ); 
nor ( n749 , n746 , n748 ); 
nand ( n750 , n745 , n749 ); 
not ( n751 , n414 ); 
nand ( n752 , n750 , n751 ); 
nor ( n753 , n752 , n358 , n416 ); 
not ( n754 , n753 ); 
not ( n755 , n393 ); 
nor ( n756 , n755 , n395 ); 
nor ( n757 , n389 , n391 ); 
and ( n758 , n756 , n757 ); 
not ( n759 , n394 ); 
nand ( n760 , n759 , n386 ); 
nand ( n761 , n758 , n760 ); 
not ( n762 , n761 ); 
nor ( n763 , n385 , n400 ); 
not ( n764 , n387 ); 
nand ( n765 , n763 , n764 ); 
not ( n766 , n765 ); 
not ( n767 , n766 ); 
not ( n768 , n767 ); 
nand ( n769 , n762 , n768 ); 
not ( n770 , n758 ); 
not ( n771 , n770 ); 
nor ( n772 , n398 , n406 ); 
nand ( n773 , n772 , n403 ); 
not ( n774 , n773 ); 
not ( n775 , n401 ); 
nand ( n776 , n774 , n775 ); 
not ( n777 , n776 ); 
nand ( n778 , n771 , n777 ); 
nand ( n779 , n769 , n778 ); 
not ( n780 , n779 ); 
or ( n781 , n754 , n780 ); 
not ( n782 , n416 ); 
not ( n783 , n782 ); 
nand ( n784 , n358 , n414 ); 
nand ( n785 , n752 , n784 ); 
not ( n786 , n785 ); 
or ( n787 , n783 , n786 ); 
not ( n788 , n311 ); 
not ( n789 , n417 ); 
not ( n790 , n789 ); 
or ( n791 , n788 , n790 ); 
not ( n792 , n311 ); 
nand ( n793 , n792 , n417 ); 
nand ( n794 , n791 , n793 ); 
not ( n795 , n794 ); 
nor ( n796 , n795 , n402 ); 
and ( n797 , n399 , n24 ); 
not ( n798 , n399 ); 
and ( n799 , n798 , n64 ); 
nor ( n800 , n797 , n799 ); 
or ( n801 , n402 , n800 ); 
nand ( n802 , n372 , n402 ); 
nand ( n803 , n801 , n802 ); 
nor ( n804 , n796 , n803 ); 
not ( n805 , n804 ); 
not ( n806 , n407 ); 
nand ( n807 , n805 , n806 ); 
nand ( n808 , n787 , n807 ); 
nand ( n809 , n808 , n762 , n406 ); 
nand ( n810 , n781 , n809 ); 
not ( n811 , n810 ); 
nor ( n812 , n397 , n390 , n405 ); 
buf ( n813 , n812 ); 
buf ( n814 , n813 ); 
not ( n815 , n814 ); 
nand ( n816 , n265 , n281 ); 
not ( n817 , n816 ); 
not ( n818 , n412 ); 
nand ( n819 , n817 , n818 ); 
not ( n820 , n819 ); 
not ( n821 , n410 ); 
nand ( n822 , n820 , n821 ); 
nor ( n823 , n392 , n815 , n822 ); 
not ( n824 , n823 ); 
or ( n825 , n811 , n824 ); 
nand ( n826 , n729 , n391 ); 
not ( n827 , n826 ); 
not ( n828 , n728 ); 
or ( n829 , n827 , n828 ); 
not ( n830 , n716 ); 
nand ( n831 , n829 , n830 ); 
nand ( n832 , n390 , n394 ); 
not ( n833 , n832 ); 
nand ( n834 , n833 , n395 ); 
and ( n835 , n831 , n834 ); 
not ( n836 , n388 ); 
or ( n837 , n836 , n816 ); 
nor ( n838 , n835 , n837 ); 
nor ( n839 , n358 , n372 ); 
buf ( n840 , n839 ); 
not ( n841 , n24 ); 
nand ( n842 , n841 , n64 ); 
not ( n843 , n842 ); 
nand ( n844 , n840 , n843 , n311 ); 
not ( n845 , n844 ); 
not ( n846 , n389 ); 
not ( n847 , n846 ); 
nand ( n848 , n373 , n715 ); 
not ( n849 , n848 ); 
not ( n850 , n849 ); 
or ( n851 , n847 , n850 ); 
nor ( n852 , n373 , n391 ); 
and ( n853 , n830 , n852 ); 
nor ( n854 , n853 , n833 ); 
nand ( n855 , n851 , n854 ); 
nand ( n856 , n845 , n855 , n393 ); 
not ( n857 , n391 ); 
not ( n858 , n857 ); 
not ( n859 , n725 ); 
or ( n860 , n858 , n859 ); 
nand ( n861 , n722 , n846 ); 
nand ( n862 , n860 , n861 ); 
nor ( n863 , n398 , n403 ); 
and ( n864 , n862 , n863 ); 
nor ( n865 , n398 , n401 ); 
not ( n866 , n865 ); 
or ( n867 , n736 , n866 ); 
nand ( n868 , n867 , n766 ); 
not ( n869 , n866 ); 
nand ( n870 , n869 , n395 ); 
nand ( n871 , n868 , n870 ); 
nor ( n872 , n864 , n871 ); 
and ( n873 , n856 , n872 ); 
nor ( n874 , n873 , n837 ); 
nor ( n875 , n838 , n874 ); 
nand ( n876 , n825 , n875 ); 
nor ( n877 , n739 , n876 ); 
not ( n878 , n774 ); 
nor ( n879 , n729 , n395 ); 
not ( n880 , n879 ); 
nor ( n881 , t_0 , n767 ); 
not ( n882 , n406 ); 
nand ( n883 , n882 , n398 ); 
nor ( n884 , n883 , n401 ); 
nand ( n885 , n765 , n884 ); 
not ( n886 , n403 ); 
not ( n887 , n886 ); 
nor ( n888 , n44 , n344 ); 
not ( n889 , n888 ); 
or ( n890 , n887 , n889 ); 
nand ( n891 , n44 , n403 ); 
nand ( n892 , n890 , n891 ); 
not ( n893 , n716 ); 
or ( n894 , n885 , n892 , n893 ); 
not ( n895 , n390 ); 
not ( n896 , n389 ); 
or ( n897 , n895 , n896 ); 
or ( n898 , n735 , n759 ); 
nand ( n899 , n897 , n898 ); 
nand ( n900 , n899 , n406 ); 
nor ( n901 , n397 , n405 ); 
not ( n902 , n901 ); 
not ( n903 , n902 ); 
nand ( n904 , n894 , n900 , n903 ); 
nor ( n905 , n881 , n904 ); 
nand ( n906 , n726 , n723 ); 
not ( n907 , n906 ); 
and ( n908 , n730 , n727 ); 
nand ( n909 , n907 , n908 ); 
not ( n910 , n24 ); 
nor ( n911 , n910 , n64 ); 
not ( n912 , n911 ); 
nand ( n913 , n912 , n842 , n358 ); 
not ( n914 , n913 ); 
nor ( n915 , n398 , n401 ); 
not ( n916 , n915 ); 
or ( n917 , n914 , n916 ); 
not ( n918 , n398 ); 
or ( n919 , n717 , n918 ); 
nand ( n920 , n917 , n919 ); 
nand ( n921 , n909 , n920 ); 
not ( n922 , n816 ); 
nor ( n923 , n922 , n913 ); 
and ( n924 , n398 , n401 ); 
nor ( n925 , n924 , n406 ); 
or ( n926 , n923 , n925 ); 
and ( n927 , n882 , n403 ); 
nand ( n928 , n927 , n401 , n918 , n888 ); 
or ( n929 , n766 , n928 ); 
nand ( n930 , n926 , n929 ); 
buf ( n931 , n862 ); 
nand ( n932 , n930 , n931 ); 
nand ( n933 , n905 , n921 , n932 ); 
nand ( n934 , n933 , n388 ); 
not ( n935 , n863 ); 
nor ( n936 , n836 , n935 ); 
nand ( n937 , n732 , n936 ); 
or ( n938 , n728 , n882 ); 
nor ( n939 , n888 , n403 ); 
not ( n940 , n939 ); 
nand ( n941 , n401 , n888 ); 
nand ( n942 , n940 , n941 ); 
not ( n943 , n942 ); 
nand ( n944 , n943 , n925 ); 
nor ( n945 , n389 , n393 ); 
nand ( n946 , n944 , n945 ); 
nand ( n947 , n938 , n946 ); 
and ( n948 , n947 , n388 ); 
nand ( n949 , n388 , n715 ); 
nor ( n950 , n949 , n817 ); 
not ( n951 , n950 ); 
not ( n952 , n951 ); 
nor ( n953 , n389 , n391 ); 
nor ( n954 , n393 , n395 ); 
nand ( n955 , n953 , n954 ); 
not ( n956 , n955 ); 
nand ( n957 , n24 , n64 ); 
nand ( n958 , n956 , n957 ); 
not ( n959 , n958 ); 
and ( n960 , n952 , n959 ); 
and ( n961 , n893 , n945 ); 
and ( n962 , n833 , n729 ); 
nor ( n963 , n961 , n962 ); 
nor ( n964 , n963 , n837 ); 
not ( n965 , n839 ); 
not ( n966 , n311 ); 
not ( n967 , n966 ); 
and ( n968 , n965 , n967 ); 
and ( n969 , n966 , n839 ); 
nor ( n970 , n968 , n969 ); 
or ( n971 , n970 , n24 ); 
not ( n972 , n64 ); 
nand ( n973 , n972 , n311 ); 
nand ( n974 , n971 , n973 , n329 ); 
and ( n975 , n964 , n974 ); 
nor ( n976 , n960 , n975 ); 
nand ( n977 , n765 , n388 ); 
not ( n978 , n395 ); 
nand ( n979 , n978 , n846 , n393 ); 
or ( n980 , n977 , n979 ); 
nand ( n981 , n980 , n837 ); 
nand ( n982 , n716 , n865 ); 
nand ( n983 , n982 , n832 ); 
nand ( n984 , n981 , n983 , n391 ); 
or ( n985 , n977 , n832 , n24 ); 
not ( n986 , n911 ); 
not ( n987 , n986 ); 
nor ( n988 , n836 , n832 ); 
nand ( n989 , n987 , n988 ); 
nand ( n990 , n985 , n989 ); 
nor ( n991 , n393 , n395 ); 
and ( n992 , n991 , n857 ); 
not ( n993 , n816 ); 
buf ( n994 , n993 ); 
not ( n995 , n994 ); 
nand ( n996 , n990 , n992 , n995 ); 
nand ( n997 , n976 , n984 , n996 ); 
nor ( n998 , n948 , n997 ); 
nand ( n999 , n857 , n389 ); 
not ( n1000 , n999 ); 
not ( n1001 , n395 ); 
nand ( n1002 , n1001 , n393 ); 
not ( n1003 , n373 ); 
nor ( n1004 , n1002 , n1003 ); 
nand ( n1005 , n1000 , n1004 ); 
nand ( n1006 , n394 , n718 ); 
or ( n1007 , n1005 , n994 , n1006 ); 
not ( n1008 , n888 ); 
buf ( n1009 , n1008 ); 
or ( n1010 , n728 , n1009 ); 
nand ( n1011 , n1007 , n1010 ); 
nand ( n1012 , n1011 , n714 ); 
nand ( n1013 , n934 , n937 , n998 , n1012 ); 
not ( n1014 , n403 ); 
nor ( n1015 , n1014 , n398 , n406 ); 
nand ( n1016 , n765 , n1015 ); 
not ( n1017 , n1016 ); 
nand ( n1018 , n718 , n44 ); 
not ( n1019 , n1018 ); 
buf ( n1020 , n1019 ); 
nand ( n1021 , n1017 , n1020 ); 
not ( n1022 , n770 ); 
nand ( n1023 , n1022 , n401 ); 
nor ( n1024 , n1021 , n1023 ); 
and ( n1025 , n1024 , n844 ); 
not ( n1026 , n415 ); 
nor ( n1027 , n1026 , n416 ); 
not ( n1028 , n1027 ); 
not ( n1029 , n407 ); 
nand ( n1030 , n1029 , n404 ); 
and ( n1031 , n1028 , n1030 ); 
nor ( n1032 , n1025 , n1031 ); 
nor ( n1033 , n388 , n410 ); 
and ( n1034 , n812 , n1033 ); 
not ( n1035 , n392 ); 
nand ( n1036 , n1034 , n1035 ); 
not ( n1037 , n1036 ); 
nand ( n1038 , n1037 , n820 ); 
not ( n1039 , n1038 ); 
and ( n1040 , n1032 , n1039 ); 
not ( n1041 , n714 ); 
nor ( n1042 , n1016 , n830 ); 
not ( n1043 , n1042 ); 
nand ( n1044 , n44 , n344 ); 
or ( n1045 , n1043 , n1044 ); 
or ( n1046 , n918 , n727 ); 
nand ( n1047 , n1045 , n1046 ); 
not ( n1048 , n1047 ); 
or ( n1049 , n1041 , n1048 ); 
or ( n1050 , n942 , n915 ); 
nand ( n1051 , n1050 , n862 ); 
not ( n1052 , n1051 ); 
not ( n1053 , n767 ); 
or ( n1054 , n1052 , n1053 ); 
nor ( n1055 , n914 , n836 ); 
nand ( n1056 , n1054 , n1055 ); 
nand ( n1057 , n1049 , n1056 ); 
nor ( n1058 , n1040 , n1057 ); 
nand ( n1059 , n956 , n329 ); 
nand ( n1060 , n778 , n1059 ); 
not ( n1061 , n1060 ); 
not ( n1062 , n1020 ); 
not ( n1063 , n398 ); 
nand ( n1064 , n1063 , n403 ); 
not ( n1065 , n1064 ); 
not ( n1066 , n1065 ); 
or ( n1067 , n1062 , n1066 ); 
nand ( n1068 , n1067 , n762 ); 
nand ( n1069 , n386 , n394 ); 
nand ( n1070 , n777 , n1069 ); 
nand ( n1071 , n1068 , n1070 ); 
not ( n1072 , n1071 ); 
nand ( n1073 , n1061 , n1072 , n769 ); 
nor ( n1074 , n1038 , n807 ); 
nand ( n1075 , n1073 , n1074 ); 
not ( n1076 , n977 ); 
not ( n1077 , n373 ); 
not ( n1078 , n991 ); 
or ( n1079 , n1077 , n1078 ); 
nor ( n1080 , n1002 , n373 ); 
nor ( n1081 , n722 , n395 ); 
nor ( n1082 , n1080 , n1081 ); 
nand ( n1083 , n1079 , n1082 ); 
and ( n1084 , n1083 , n830 ); 
and ( n1085 , n983 , n727 ); 
nor ( n1086 , n1084 , n1085 ); 
or ( n1087 , n1086 , n999 ); 
not ( n1088 , n723 ); 
not ( n1089 , n979 ); 
nand ( n1090 , n1088 , n1089 ); 
or ( n1091 , n1090 , n717 ); 
nand ( n1092 , n1087 , n1091 ); 
nand ( n1093 , n1076 , n1092 ); 
nand ( n1094 , n1058 , n1075 , n1093 ); 
nor ( n1095 , n1013 , n1094 ); 
not ( n1096 , n785 ); 
and ( n1097 , n1034 , n782 ); 
not ( n1098 , n1097 ); 
nor ( n1099 , n1098 , n392 ); 
nand ( n1100 , n1099 , n820 ); 
nor ( n1101 , n1096 , n1100 ); 
and ( n1102 , n1101 , n1071 ); 
not ( n1103 , n1059 ); 
and ( n1104 , n1101 , n1103 ); 
nor ( n1105 , n1102 , n1104 ); 
not ( n1106 , n358 ); 
not ( n1107 , n750 ); 
or ( n1108 , n1106 , n1107 ); 
not ( n1109 , n784 ); 
not ( n1110 , n1109 ); 
nand ( n1111 , n1108 , n1110 ); 
and ( n1112 , n779 , n1111 ); 
nor ( n1113 , n761 , n844 ); 
not ( n1114 , n409 ); 
nand ( n1115 , n751 , n1114 ); 
not ( n1116 , n1115 ); 
nor ( n1117 , n413 , n414 ); 
nor ( n1118 , n1116 , n1117 ); 
not ( n1119 , n1118 ); 
and ( n1120 , n1113 , n1119 ); 
nor ( n1121 , n1112 , n1120 ); 
not ( n1122 , n1121 ); 
not ( n1123 , n1100 ); 
and ( n1124 , n1122 , n1123 ); 
nor ( n1125 , n402 , n407 ); 
nand ( n1126 , n399 , n417 ); 
nand ( n1127 , n1113 , n1039 , n1125 , n1126 ); 
not ( n1128 , n344 ); 
nor ( n1129 , n1016 , n775 ); 
not ( n1130 , n1129 ); 
or ( n1131 , n1128 , n1130 ); 
buf ( n1132 , n885 ); 
nand ( n1133 , n1131 , n1132 ); 
and ( n1134 , n988 , n1133 ); 
and ( n1135 , n735 , n727 ); 
and ( n1136 , n950 , n1135 ); 
nor ( n1137 , n391 , n395 ); 
not ( n1138 , n1137 ); 
nor ( n1139 , n1138 , n993 ); 
and ( n1140 , n1139 , n988 ); 
nor ( n1141 , n1136 , n1140 ); 
nor ( n1142 , n842 , n311 ); 
nand ( n1143 , n1142 , n840 ); 
or ( n1144 , n1141 , n1143 ); 
and ( n1145 , n942 , n899 ); 
and ( n1146 , n956 , n915 ); 
nor ( n1147 , n1145 , n1146 ); 
or ( n1148 , n1147 , n836 ); 
nand ( n1149 , n1144 , n1148 ); 
nor ( n1150 , n1134 , n1149 ); 
not ( n1151 , n931 ); 
nor ( n1152 , n1151 , n949 ); 
and ( n1153 , n1133 , n1152 ); 
not ( n1154 , n1000 ); 
nor ( n1155 , n359 , n373 ); 
nand ( n1156 , n954 , n1155 ); 
nand ( n1157 , n879 , n373 ); 
nand ( n1158 , n1156 , n1157 ); 
not ( n1159 , n1158 ); 
or ( n1160 , n1154 , n1159 ); 
not ( n1161 , n395 ); 
nand ( n1162 , n1161 , n846 , n393 ); 
not ( n1163 , n1162 ); 
buf ( n1164 , n725 ); 
nand ( n1165 , n1163 , n1164 , n391 ); 
nand ( n1166 , n1160 , n1165 ); 
not ( n1167 , n977 ); 
and ( n1168 , n1166 , n1167 , n390 ); 
nor ( n1169 , n1153 , n1168 ); 
nand ( n1170 , n1127 , n1150 , n1169 ); 
nor ( n1171 , n1124 , n1170 ); 
nand ( n1172 , n877 , n1095 , n1105 , n1171 ); 
not ( n1173 , n265 ); 
nor ( n1174 , n1173 , n281 ); 
nand ( n1175 , n393 , n1155 ); 
not ( n1176 , n1175 ); 
not ( n1177 , n1176 ); 
not ( n1178 , n717 ); 
not ( n1179 , n1178 ); 
or ( n1180 , n1177 , n1179 ); 
not ( n1181 , n1178 ); 
not ( n1182 , n862 ); 
or ( n1183 , n1181 , n1182 ); 
not ( n1184 , n390 ); 
not ( n1185 , n394 ); 
or ( n1186 , n1184 , n1185 ); 
nand ( n1187 , n1186 , n388 ); 
not ( n1188 , n1187 ); 
nand ( n1189 , n1183 , n1188 ); 
not ( n1190 , n1189 ); 
nand ( n1191 , n1180 , n1190 ); 
and ( n1192 , n1174 , n1191 ); 
not ( n1193 , n717 ); 
not ( n1194 , n44 ); 
nand ( n1195 , n1194 , n344 ); 
and ( n1196 , n1195 , n1018 ); 
not ( n1197 , n1196 ); 
or ( n1198 , n1193 , n1197 ); 
or ( n1199 , n1175 , n1009 ); 
nand ( n1200 , n1198 , n1199 ); 
nor ( n1201 , n1192 , n1200 ); 
not ( n1202 , n1201 ); 
and ( n1203 , n392 , n401 ); 
nand ( n1204 , n1017 , n1203 ); 
not ( n1205 , n1204 ); 
and ( n1206 , n1202 , n1205 ); 
and ( n1207 , n738 , n1203 ); 
nor ( n1208 , n1206 , n1207 ); 
nor ( n1209 , n1118 , n1126 ); 
not ( n1210 , n1209 ); 
not ( n1211 , n1113 ); 
or ( n1212 , n1210 , n1211 ); 
not ( n1213 , n1021 ); 
not ( n1214 , n402 ); 
nor ( n1215 , n1213 , n1214 ); 
not ( n1216 , n372 ); 
nand ( n1217 , n1216 , n758 ); 
not ( n1218 , n1217 ); 
and ( n1219 , n1218 , n760 ); 
not ( n1220 , n358 ); 
and ( n1221 , n751 , n1220 ); 
and ( n1222 , n281 , n358 ); 
nor ( n1223 , n1221 , n1222 ); 
not ( n1224 , n1223 ); 
nand ( n1225 , n1215 , n1219 , n744 , n1224 ); 
nand ( n1226 , n1212 , n1225 ); 
not ( n1227 , n762 ); 
not ( n1228 , n1016 ); 
nand ( n1229 , n1228 , n1020 ); 
not ( n1230 , n1229 ); 
or ( n1231 , n1227 , n1230 ); 
nand ( n1232 , n1231 , n1070 ); 
not ( n1233 , n1232 ); 
and ( n1234 , n800 , n1214 ); 
not ( n1235 , n1234 ); 
nor ( n1236 , n311 , n417 ); 
and ( n1237 , n409 , n1236 ); 
not ( n1238 , n409 ); 
nand ( n1239 , n311 , n417 ); 
not ( n1240 , n1239 ); 
and ( n1241 , n1238 , n1240 ); 
nor ( n1242 , n1237 , n1241 ); 
nor ( n1243 , n1235 , n1242 , n1223 ); 
not ( n1244 , n1243 ); 
or ( n1245 , n1233 , n1244 ); 
not ( n1246 , n751 ); 
not ( n1247 , n744 ); 
or ( n1248 , n1246 , n1247 ); 
and ( n1249 , n1117 , n64 ); 
nor ( n1250 , n1249 , n1109 ); 
nand ( n1251 , n1248 , n1250 ); 
nand ( n1252 , n1218 , n777 , n1251 , n402 ); 
nand ( n1253 , n1245 , n1252 ); 
or ( n1254 , n1226 , n1253 ); 
and ( n1255 , n1097 , n265 ); 
not ( n1256 , n404 ); 
and ( n1257 , n1255 , n1256 ); 
nand ( n1258 , n1254 , n1257 ); 
nand ( n1259 , n1208 , n1258 ); 
not ( n1260 , n265 ); 
or ( n1261 , n717 , n1260 ); 
nand ( n1262 , n1261 , n1009 ); 
and ( n1263 , n1203 , n1262 , n732 ); 
or ( n1264 , n1008 , n398 ); 
not ( n1265 , n939 ); 
nand ( n1266 , n1264 , n1265 ); 
and ( n1267 , n862 , n1266 ); 
nor ( n1268 , n1267 , n768 ); 
or ( n1269 , n1268 , n923 , n1035 ); 
not ( n1270 , n730 ); 
not ( n1271 , n723 ); 
or ( n1272 , n1270 , n1271 ); 
nand ( n1273 , n1272 , n406 ); 
not ( n1274 , n730 ); 
nand ( n1275 , n1274 , n886 , n44 ); 
and ( n1276 , n1273 , n1275 ); 
or ( n1277 , n1276 , n1035 ); 
nand ( n1278 , n1269 , n1277 ); 
nor ( n1279 , n1263 , n1278 ); 
not ( n1280 , n1255 ); 
not ( n1281 , n1256 ); 
nor ( n1282 , n1214 , n372 ); 
not ( n1283 , n1282 ); 
or ( n1284 , n1281 , n1283 ); 
nand ( n1285 , n1284 , n806 ); 
nand ( n1286 , n1214 , n399 ); 
nor ( n1287 , n1286 , n404 , n417 ); 
or ( n1288 , n1285 , n1287 ); 
not ( n1289 , n1116 ); 
not ( n1290 , n413 ); 
or ( n1291 , n1289 , n1290 ); 
nand ( n1292 , n1288 , n1291 ); 
nor ( n1293 , n761 , n1292 ); 
not ( n1294 , n1293 ); 
or ( n1295 , n1280 , n1294 ); 
and ( n1296 , n392 , n1189 ); 
not ( n1297 , n1034 ); 
and ( n1298 , n1027 , n1030 ); 
nor ( n1299 , n1298 , n412 ); 
nor ( n1300 , n1297 , n1299 ); 
nor ( n1301 , n1296 , n1300 ); 
or ( n1302 , n1301 , n1260 ); 
nand ( n1303 , n1295 , n1302 ); 
nand ( n1304 , n1303 , n1142 , n358 ); 
not ( n1305 , n899 ); 
not ( n1306 , n945 ); 
nand ( n1307 , n1003 , n393 , n389 ); 
nand ( n1308 , n1306 , n1307 ); 
not ( n1309 , n1308 ); 
and ( n1310 , n728 , n1305 , n1309 ); 
nor ( n1311 , n1310 , n935 ); 
nand ( n1312 , n857 , n1080 ); 
not ( n1313 , n359 ); 
nand ( n1314 , n1313 , n1089 ); 
and ( n1315 , n1312 , n1314 ); 
nor ( n1316 , n1315 , n1016 , n401 ); 
or ( n1317 , n1311 , n1316 ); 
nand ( n1318 , n1317 , n392 ); 
nand ( n1319 , n762 , n1021 ); 
or ( n1320 , n1319 , n806 ); 
not ( n1321 , n1285 ); 
or ( n1322 , n1070 , n1321 ); 
nand ( n1323 , n1320 , n1322 ); 
nand ( n1324 , n1323 , n1255 , n750 , n1224 ); 
nand ( n1325 , n1279 , n1304 , n1318 , n1324 ); 
nor ( n1326 , n1259 , n1325 ); 
and ( n1327 , n1219 , n1215 ); 
nor ( n1328 , n842 , n413 ); 
and ( n1329 , n1327 , n1328 ); 
not ( n1330 , n399 ); 
nand ( n1331 , n911 , n1330 ); 
not ( n1332 , n1331 ); 
nand ( n1333 , n1332 , n1219 ); 
nand ( n1334 , n795 , n413 ); 
nor ( n1335 , n1333 , n1334 ); 
nor ( n1336 , n1329 , n1335 ); 
or ( n1337 , n1232 , n1060 ); 
nor ( n1338 , n1334 , n1331 , n402 ); 
nor ( n1339 , n794 , n1286 ); 
and ( n1340 , n1339 , n1328 ); 
or ( n1341 , n1338 , n1340 ); 
nand ( n1342 , n1337 , n1341 ); 
and ( n1343 , n1336 , n1342 ); 
nand ( n1344 , n1257 , n751 ); 
nor ( n1345 , n1343 , n1344 ); 
nor ( n1346 , n1260 , n281 ); 
nand ( n1347 , n1034 , n1346 ); 
not ( n1348 , n1347 ); 
nand ( n1349 , n765 , n927 ); 
not ( n1350 , n1349 ); 
and ( n1351 , n1348 , n1350 ); 
and ( n1352 , n1042 , n392 ); 
nor ( n1353 , n1351 , n1352 ); 
or ( n1354 , n1089 , n1137 ); 
nand ( n1355 , n1354 , n775 ); 
or ( n1356 , n1353 , n1355 ); 
not ( n1357 , n716 ); 
nor ( n1358 , n1357 , n1187 ); 
or ( n1359 , n1358 , n958 ); 
nor ( n1360 , n1308 , n395 ); 
or ( n1361 , n1360 , n925 ); 
nand ( n1362 , n1359 , n1361 ); 
and ( n1363 , n1362 , n392 ); 
nand ( n1364 , n992 , n869 ); 
not ( n1365 , n1188 ); 
not ( n1366 , n848 ); 
or ( n1367 , n1365 , n1366 ); 
nor ( n1368 , n1162 , n857 ); 
nand ( n1369 , n1367 , n1368 ); 
and ( n1370 , n1364 , n1369 ); 
nor ( n1371 , n766 , n1035 ); 
nand ( n1372 , n1371 , n359 ); 
nor ( n1373 , n1370 , n1372 ); 
nor ( n1374 , n1363 , n1373 ); 
nand ( n1375 , n1356 , n1374 ); 
nand ( n1376 , n1166 , n1371 , n390 ); 
not ( n1377 , n1006 ); 
nand ( n1378 , n1377 , n1166 , n1203 ); 
nand ( n1379 , n1376 , n1378 ); 
nand ( n1380 , n1300 , n994 ); 
or ( n1381 , n1024 , n1380 ); 
or ( n1382 , n970 , n842 , n265 ); 
or ( n1383 , n1382 , n1358 ); 
nand ( n1384 , n1383 , n776 ); 
nand ( n1385 , n1384 , n1135 , n392 ); 
nand ( n1386 , n1381 , n1385 ); 
nor ( n1387 , n1375 , n1379 , n1386 ); 
not ( n1388 , n1234 ); 
or ( n1389 , n1388 , n404 , n794 ); 
nand ( n1390 , n1389 , n1321 ); 
and ( n1391 , n1097 , n1390 , n994 , n1109 ); 
and ( n1392 , n1391 , n1232 ); 
and ( n1393 , n833 , n727 , n373 ); 
nand ( n1394 , n848 , n388 ); 
and ( n1395 , n1394 , n991 ); 
nor ( n1396 , n1393 , n1395 ); 
or ( n1397 , n1396 , n999 , n359 ); 
or ( n1398 , n1005 , n388 ); 
nand ( n1399 , n1397 , n1398 ); 
and ( n1400 , n1399 , n1371 ); 
nor ( n1401 , n1392 , n1400 ); 
or ( n1402 , n778 , n806 ); 
or ( n1403 , n1321 , n1059 ); 
nand ( n1404 , n1402 , n1403 ); 
and ( n1405 , n1255 , n1404 , n785 ); 
not ( n1406 , n1129 ); 
and ( n1407 , n1132 , n914 ); 
nand ( n1408 , n777 , n1135 ); 
buf ( n1409 , n770 ); 
nand ( n1410 , n776 , n1409 ); 
nand ( n1411 , n1406 , n1407 , n1408 , n1410 ); 
not ( n1412 , n1347 ); 
and ( n1413 , n1411 , n1412 ); 
nor ( n1414 , n1405 , n1413 ); 
nand ( n1415 , n1387 , n1401 , n1414 ); 
nor ( n1416 , n1345 , n1415 ); 
not ( n1417 , n1234 ); 
not ( n1418 , n1060 ); 
or ( n1419 , n1417 , n1418 ); 
nand ( n1420 , n1419 , n1333 ); 
and ( n1421 , n1420 , n1257 ); 
not ( n1422 , n1236 ); 
not ( n1423 , n409 ); 
nor ( n1424 , n1423 , n414 ); 
not ( n1425 , n1424 ); 
or ( n1426 , n1422 , n1425 ); 
or ( n1427 , n794 , n1110 ); 
or ( n1428 , n1239 , n1289 ); 
nand ( n1429 , n1426 , n1427 , n1428 ); 
and ( n1430 , n1421 , n1429 ); 
nand ( n1431 , n840 , n64 , n311 ); 
or ( n1432 , n1431 , n1118 ); 
nand ( n1433 , n745 , n1290 ); 
nand ( n1434 , n1433 , n840 , n751 , n24 ); 
nand ( n1435 , n1432 , n1434 ); 
and ( n1436 , n762 , n1435 ); 
and ( n1437 , n358 , n1433 ); 
nor ( n1438 , n1437 , n1109 ); 
or ( n1439 , n1438 , n986 ); 
or ( n1440 , n1223 , n957 ); 
nand ( n1441 , n1439 , n1440 ); 
and ( n1442 , n1219 , n1441 ); 
nor ( n1443 , n1436 , n1442 ); 
not ( n1444 , n1255 ); 
and ( n1445 , n1256 , n402 ); 
nor ( n1446 , n1445 , n407 ); 
or ( n1447 , n1443 , n1444 , n1446 ); 
not ( n1448 , n372 ); 
and ( n1449 , n994 , n1448 , n24 ); 
nor ( n1450 , n1431 , n1260 ); 
nor ( n1451 , n1449 , n1450 ); 
or ( n1452 , n1301 , n1451 ); 
nand ( n1453 , n1447 , n1452 ); 
nor ( n1454 , n1430 , n1453 ); 
and ( n1455 , n905 , n921 , n932 ); 
not ( n1456 , n1455 ); 
or ( n1457 , n1309 , n716 ); 
not ( n1458 , n1409 ); 
or ( n1459 , n1458 , n1188 ); 
and ( n1460 , n906 , n915 ); 
nand ( n1461 , n870 , n982 ); 
nor ( n1462 , n1460 , n1461 ); 
nand ( n1463 , n1457 , n1459 , n1462 ); 
and ( n1464 , n1463 , n994 ); 
and ( n1465 , n1133 , n1191 ); 
nor ( n1466 , n1464 , n1465 ); 
not ( n1467 , n1466 ); 
or ( n1468 , n1456 , n1467 ); 
nand ( n1469 , n1468 , n392 ); 
nand ( n1470 , n1326 , n1416 , n1454 , n1469 ); 
not ( n1471 , n1006 ); 
and ( n1472 , n1166 , n1471 ); 
not ( n1473 , n401 ); 
nor ( n1474 , n1473 , n390 ); 
and ( n1475 , n1472 , n1474 ); 
nor ( n1476 , n1475 , n836 ); 
not ( n1477 , n1476 ); 
not ( n1478 , n400 ); 
nor ( n1479 , n1478 , n387 ); 
and ( n1480 , n1477 , n1479 ); 
nor ( n1481 , n775 , n406 ); 
nand ( n1482 , n1004 , n1481 ); 
not ( n1483 , n401 ); 
not ( n1484 , n878 ); 
or ( n1485 , n1483 , n1484 ); 
not ( n1486 , n1156 ); 
nand ( n1487 , n1485 , n1486 ); 
nand ( n1488 , n1482 , n1487 ); 
and ( n1489 , n813 , n388 ); 
nor ( n1490 , n846 , n394 ); 
nand ( n1491 , n1488 , n1489 , n1490 ); 
nand ( n1492 , n774 , n401 ); 
not ( n1493 , n1492 ); 
not ( n1494 , n397 ); 
not ( n1495 , n405 ); 
nand ( n1496 , n1494 , n1495 ); 
nor ( n1497 , n999 , n1496 ); 
not ( n1498 , n1195 ); 
nand ( n1499 , n1158 , n1493 , n1497 , n1498 ); 
and ( n1500 , n391 , n394 ); 
or ( n1501 , n892 , n918 ); 
or ( n1502 , n1498 , n775 ); 
nand ( n1503 , n1501 , n1502 ); 
nand ( n1504 , n1489 , n1500 , n1503 ); 
nand ( n1505 , n1491 , n1499 , n1504 ); 
nand ( n1506 , n1019 , n389 ); 
nor ( n1507 , n1157 , n1506 ); 
not ( n1508 , n1507 ); 
not ( n1509 , n1493 ); 
or ( n1510 , n1508 , n1509 ); 
nand ( n1511 , n1164 , n1089 ); 
and ( n1512 , n759 , n391 ); 
nand ( n1513 , n1511 , n1512 ); 
nand ( n1514 , n1510 , n1513 ); 
nand ( n1515 , n1514 , n1489 ); 
or ( n1516 , n863 , n882 ); 
or ( n1517 , n775 , n403 ); 
nand ( n1518 , n1516 , n1517 ); 
nand ( n1519 , n1489 , n1518 , n1500 ); 
and ( n1520 , n1486 , n1000 ); 
and ( n1521 , n892 , n884 , n901 ); 
nand ( n1522 , n1520 , n1521 ); 
nand ( n1523 , n1515 , n1519 , n1522 ); 
nor ( n1524 , n1505 , n1523 ); 
and ( n1525 , n385 , n387 ); 
nand ( n1526 , n1525 , n1478 ); 
or ( n1527 , n1524 , n1526 ); 
and ( n1528 , n1497 , n836 ); 
not ( n1529 , n1528 ); 
not ( n1530 , n775 ); 
not ( n1531 , n398 ); 
or ( n1532 , n1530 , n1531 ); 
nand ( n1533 , n1532 , n1492 ); 
not ( n1534 , n1533 ); 
not ( n1535 , n1486 ); 
or ( n1536 , n1534 , n1535 ); 
nand ( n1537 , n1536 , n1482 ); 
not ( n1538 , n1537 ); 
or ( n1539 , n1529 , n1538 ); 
nand ( n1540 , n775 , n406 ); 
not ( n1541 , n1540 ); 
nand ( n1542 , n1541 , n991 , n935 ); 
nand ( n1543 , n879 , n1064 , n1481 ); 
nand ( n1544 , n1542 , n1543 ); 
nand ( n1545 , n1528 , n1544 ); 
nand ( n1546 , n1539 , n1545 ); 
and ( n1547 , n1546 , n1525 ); 
nand ( n1548 , n1479 , n397 ); 
and ( n1549 , n392 , n414 ); 
not ( n1550 , n392 ); 
and ( n1551 , n1550 , n402 ); 
or ( n1552 , n1549 , n1551 ); 
nor ( n1553 , n1548 , n1552 ); 
nor ( n1554 , n1547 , n1553 ); 
nand ( n1555 , n1527 , n1554 ); 
nor ( n1556 , n1480 , n1555 ); 
not ( n1557 , n1020 ); 
not ( n1558 , n1482 ); 
not ( n1559 , n1558 ); 
or ( n1560 , n1557 , n1559 ); 
not ( n1561 , n1544 ); 
nand ( n1562 , n1560 , n1561 ); 
and ( n1563 , n1562 , n1000 ); 
nor ( n1564 , n1563 , t_1 ); 
not ( n1565 , n390 ); 
nor ( n1566 , n1564 , n1565 ); 
not ( n1567 , n1566 ); 
nor ( n1568 , n999 , n832 ); 
nand ( n1569 , n1537 , n1568 ); 
and ( n1570 , n1567 , n1569 ); 
nor ( n1571 , n1570 , n405 ); 
nor ( n1572 , n1494 , n405 ); 
nand ( n1573 , n390 , n1572 ); 
not ( n1574 , n1573 ); 
or ( n1575 , n1571 , n1574 ); 
not ( n1576 , n1526 ); 
nand ( n1577 , n1575 , n1576 ); 
and ( n1578 , n729 , n373 ); 
nor ( n1579 , n1578 , n1176 ); 
not ( n1580 , n1579 ); 
not ( n1581 , n731 ); 
or ( n1582 , n1580 , n1581 ); 
nand ( n1583 , n1582 , n1193 ); 
not ( n1584 , n1583 ); 
not ( n1585 , n1525 ); 
nand ( n1586 , n1584 , n1585 , n400 ); 
and ( n1587 , n1472 , n401 ); 
nor ( n1588 , n1587 , n397 ); 
not ( n1589 , n385 ); 
nand ( n1590 , n1589 , n400 ); 
nor ( n1591 , n1588 , n1590 ); 
nand ( n1592 , n1494 , n390 ); 
not ( n1593 , n1592 ); 
not ( n1594 , n1593 ); 
not ( n1595 , n1166 ); 
or ( n1596 , n1594 , n1595 ); 
not ( n1597 , n863 ); 
not ( n1598 , n775 ); 
or ( n1599 , n1597 , n1598 ); 
nand ( n1600 , n865 , n882 ); 
nand ( n1601 , n1599 , n1600 ); 
not ( n1602 , n390 ); 
nand ( n1603 , n1602 , n394 ); 
nand ( n1604 , n1603 , n1592 ); 
and ( n1605 , n1601 , n1604 ); 
or ( n1606 , n1494 , n390 ); 
nand ( n1607 , n1606 , n1495 ); 
nor ( n1608 , n1605 , n1607 ); 
nand ( n1609 , n393 , n395 ); 
and ( n1610 , n1609 , n736 ); 
not ( n1611 , n1609 ); 
and ( n1612 , n1611 , n999 ); 
nor ( n1613 , n1610 , n1612 ); 
nand ( n1614 , n1613 , n893 ); 
nand ( n1615 , n1187 , n1494 ); 
and ( n1616 , n1608 , n1614 , n1615 ); 
nand ( n1617 , n1596 , n1616 ); 
not ( n1618 , n1617 ); 
not ( n1619 , n1008 ); 
not ( n1620 , n886 ); 
and ( n1621 , n1619 , n1620 ); 
or ( n1622 , n1195 , n401 ); 
or ( n1623 , n1044 , n775 ); 
nand ( n1624 , n1622 , n1623 ); 
nor ( n1625 , n1621 , n1624 ); 
and ( n1626 , n943 , n1625 , n925 ); 
not ( n1627 , n387 ); 
and ( n1628 , n1604 , n1627 ); 
and ( n1629 , n716 , n1589 ); 
nor ( n1630 , n1628 , n1629 ); 
or ( n1631 , n1626 , n1630 ); 
not ( n1632 , n1593 ); 
nor ( n1633 , n1632 , n1613 ); 
nand ( n1634 , n1633 , n1525 ); 
nand ( n1635 , n1631 , n1634 ); 
not ( n1636 , n1635 ); 
and ( n1637 , n1618 , n1636 ); 
nor ( n1638 , n1637 , n1478 ); 
nor ( n1639 , n1591 , n1638 ); 
nand ( n1640 , n1556 , n1577 , n1586 , n1639 ); 
not ( n1641 , n1626 ); 
and ( n1642 , n1641 , n1604 ); 
nor ( n1643 , n1552 , n400 ); 
not ( n1644 , n1643 ); 
and ( n1645 , n1644 , n397 ); 
nor ( n1646 , n1642 , n1645 ); 
nand ( n1647 , n1476 , n1583 , n1646 ); 
nor ( n1648 , n1627 , n385 ); 
nand ( n1649 , n1647 , n1648 ); 
buf ( n1650 , n903 ); 
not ( n1651 , n1650 ); 
not ( n1652 , n1566 ); 
or ( n1653 , n1651 , n1652 ); 
not ( n1654 , n1497 ); 
not ( n1655 , n1654 ); 
and ( n1656 , n1537 , n1655 , n1187 ); 
not ( n1657 , n1545 ); 
nor ( n1658 , n1656 , n1657 ); 
nand ( n1659 , n1653 , n1658 ); 
and ( n1660 , n385 , n1659 ); 
not ( n1661 , n387 ); 
nand ( n1662 , n1661 , n385 ); 
or ( n1663 , n1524 , n1662 ); 
nand ( n1664 , n1617 , n387 ); 
or ( n1665 , n1573 , n1552 ); 
not ( n1666 , n388 ); 
nand ( n1667 , n1666 , n390 ); 
not ( n1668 , n1667 ); 
nand ( n1669 , n1668 , n1572 ); 
nand ( n1670 , n1665 , n1669 ); 
and ( n1671 , n1479 , n385 ); 
and ( n1672 , n1670 , n1671 ); 
nor ( n1673 , n1573 , n836 ); 
nor ( n1674 , n1662 , n400 ); 
and ( n1675 , n1673 , n1674 ); 
nor ( n1676 , n1672 , n1675 ); 
and ( n1677 , n1676 , n1634 ); 
nand ( n1678 , n1663 , n1664 , n1677 ); 
nor ( n1679 , n1660 , n1678 ); 
nand ( n1680 , n1649 , n1679 ); 
not ( n1681 , n995 ); 
nand ( n1682 , n408 , n412 ); 
not ( n1683 , n1682 ); 
and ( n1684 , n1681 , n1683 ); 
nand ( n1685 , n1218 , n914 ); 
not ( n1686 , n412 ); 
and ( n1687 , n1686 , n311 ); 
not ( n1688 , n1687 ); 
or ( n1689 , n1688 , n281 ); 
or ( n1690 , n1260 , n1682 ); 
or ( n1691 , n265 , n966 ); 
nand ( n1692 , n1689 , n1690 , n1691 ); 
and ( n1693 , n1685 , n1692 ); 
nor ( n1694 , n1684 , n1693 ); 
not ( n1695 , n1694 ); 
not ( n1696 , n1036 ); 
and ( n1697 , n1695 , n1696 ); 
nand ( n1698 , n923 , n1218 ); 
nor ( n1699 , n388 , n392 ); 
or ( n1700 , n1699 , n759 ); 
nand ( n1701 , n1700 , n832 ); 
nand ( n1702 , n1698 , n1701 ); 
nor ( n1703 , n1290 , n24 ); 
and ( n1704 , n1703 , n399 ); 
nor ( n1705 , n24 , n64 ); 
nor ( n1706 , n1704 , n1705 ); 
not ( n1707 , n1706 ); 
not ( n1708 , n372 ); 
not ( n1709 , n394 ); 
nor ( n1710 , n1709 , n410 ); 
nand ( n1711 , n1687 , n1710 , n417 ); 
nor ( n1712 , n1711 , n1425 , n402 ); 
not ( n1713 , n1712 ); 
or ( n1714 , n1708 , n1713 ); 
not ( n1715 , n1710 ); 
nor ( n1716 , n819 , n1715 ); 
nand ( n1717 , n1236 , n1256 ); 
nand ( n1718 , n1214 , n1026 ); 
nor ( n1719 , n1717 , n1115 , n1718 ); 
nand ( n1720 , n1716 , n1719 ); 
nand ( n1721 , n1714 , n1720 ); 
nand ( n1722 , n1707 , n1721 ); 
nor ( n1723 , n1331 , n413 ); 
not ( n1724 , n1723 ); 
not ( n1725 , n1712 ); 
or ( n1726 , n1724 , n1725 ); 
nor ( n1727 , n751 , n358 ); 
nand ( n1728 , n1727 , n1026 ); 
nand ( n1729 , n372 , n416 ); 
and ( n1730 , n1728 , n1729 ); 
nor ( n1731 , n1730 , n1711 ); 
nand ( n1732 , n1731 , n1234 ); 
nand ( n1733 , n1726 , n1732 ); 
not ( n1734 , n902 ); 
or ( n1735 , n1734 , n759 ); 
nor ( n1736 , n1715 , n1290 , n1126 , n372 ); 
nand ( n1737 , n1736 , n1424 , n1687 , n843 ); 
nand ( n1738 , n1735 , n1737 ); 
nor ( n1739 , n1733 , n1738 ); 
nand ( n1740 , n1702 , n1722 , n1739 ); 
nor ( n1741 , n1697 , n1740 ); 
not ( n1742 , n1135 ); 
not ( n1743 , n1600 ); 
not ( n1744 , n396 ); 
or ( n1745 , n1743 , n1744 ); 
or ( n1746 , n329 , n393 ); 
nand ( n1747 , n1745 , n1746 ); 
nor ( n1748 , n1742 , n1747 ); 
and ( n1749 , n1256 , n416 ); 
and ( n1750 , n1030 , n1026 ); 
nor ( n1751 , n1749 , n1750 ); 
or ( n1752 , n1748 , n1751 ); 
not ( n1753 , n1705 ); 
not ( n1754 , n1424 ); 
or ( n1755 , n1753 , n1754 ); 
nand ( n1756 , n800 , n416 ); 
nand ( n1757 , n1755 , n1756 ); 
nand ( n1758 , n1757 , n1240 , n1448 ); 
nand ( n1759 , n1752 , n1758 ); 
and ( n1760 , n1759 , n1716 ); 
nand ( n1761 , n1716 , n1285 , n749 ); 
nor ( n1762 , n1761 , n1289 , n311 , n415 ); 
not ( n1763 , n311 ); 
nor ( n1764 , n1761 , n1763 , n1425 ); 
nor ( n1765 , n1760 , n1762 , n1764 ); 
and ( n1766 , n814 , n1699 , n410 , n411 ); 
and ( n1767 , n1698 , n1766 ); 
or ( n1768 , n1388 , n1717 ); 
nand ( n1769 , n1768 , n1321 ); 
and ( n1770 , n1728 , n782 ); 
not ( n1771 , n1716 ); 
nor ( n1772 , n1770 , n1771 ); 
and ( n1773 , n1769 , n1772 ); 
not ( n1774 , n1720 ); 
nor ( n1775 , n399 , n64 , n413 ); 
and ( n1776 , n1774 , n1775 ); 
nor ( n1777 , n1767 , n1773 , n1776 ); 
and ( n1778 , n1741 , n1765 , n1777 ); 
nand ( n1779 , n777 , n396 ); 
not ( n1780 , n1779 ); 
nand ( n1781 , n1780 , n358 ); 
nor ( n1782 , n1100 , n1781 ); 
nand ( n1783 , n1782 , n409 ); 
not ( n1784 , n1783 ); 
not ( n1785 , n1026 ); 
nand ( n1786 , n1687 , n1220 ); 
nor ( n1787 , n1779 , n1786 ); 
not ( n1788 , n1787 ); 
or ( n1789 , n1785 , n1788 ); 
nor ( n1790 , n329 , n1688 , n955 ); 
and ( n1791 , n777 , n1790 ); 
nand ( n1792 , n1791 , n1028 ); 
nand ( n1793 , n1789 , n1792 ); 
not ( n1794 , n1036 ); 
and ( n1795 , n1793 , n1794 ); 
and ( n1796 , n1039 , n1780 , n311 , n416 ); 
nor ( n1797 , n1795 , n1796 ); 
not ( n1798 , n1797 ); 
or ( n1799 , n1784 , n1798 ); 
and ( n1800 , n806 , n1256 ); 
not ( n1801 , n1800 ); 
nor ( n1802 , n1801 , n402 , n417 ); 
nand ( n1803 , n1799 , n1802 ); 
or ( n1804 , n414 , n749 ); 
nand ( n1805 , n1804 , n1110 ); 
and ( n1806 , n1805 , n1750 ); 
not ( n1807 , n1030 ); 
nor ( n1808 , n1425 , n1807 , n311 ); 
nor ( n1809 , n1806 , n1808 ); 
or ( n1810 , n1100 , n1809 ); 
and ( n1811 , n803 , n1800 ); 
not ( n1812 , n793 ); 
and ( n1813 , n1812 , n1125 ); 
nor ( n1814 , n1811 , n1813 ); 
not ( n1815 , n1814 ); 
nand ( n1816 , n1815 , n1028 ); 
or ( n1817 , n1038 , n1816 ); 
nand ( n1818 , n1810 , n1817 ); 
or ( n1819 , n776 , n955 , n329 ); 
nand ( n1820 , n1819 , n1779 ); 
and ( n1821 , n1818 , n1820 ); 
nand ( n1822 , n1039 , n1030 , n1027 , n409 ); 
nand ( n1823 , n1039 , n1807 , n417 ); 
nand ( n1824 , n1822 , n1823 ); 
nor ( n1825 , n1821 , n1824 ); 
nor ( n1826 , n1763 , n409 ); 
not ( n1827 , n1826 ); 
not ( n1828 , n1782 ); 
or ( n1829 , n1827 , n1828 ); 
or ( n1830 , n1787 , n1791 ); 
nand ( n1831 , n1830 , n1099 , n1116 ); 
nand ( n1832 , n1829 , n1831 ); 
nand ( n1833 , n1832 , n1750 ); 
nand ( n1834 , n1778 , n1803 , n1825 , n1833 ); 
nand ( n1835 , n782 , n1026 ); 
nor ( n1836 , n1835 , n1807 ); 
and ( n1837 , n785 , n1836 ); 
buf ( n1838 , n804 ); 
nand ( n1839 , n1028 , n1800 ); 
nor ( n1840 , n1838 , n1839 ); 
nor ( n1841 , n1837 , n1840 ); 
and ( n1842 , n1135 , n329 ); 
nor ( n1843 , n1842 , n1410 ); 
or ( n1844 , n1841 , n1038 , n1843 ); 
not ( n1845 , n822 ); 
not ( n1846 , n388 ); 
and ( n1847 , n1845 , n1846 ); 
nor ( n1848 , n1667 , n392 ); 
nand ( n1849 , n281 , n1686 , n1848 ); 
nand ( n1850 , n1033 , n392 , n265 , n390 ); 
nand ( n1851 , n1849 , n1850 ); 
nor ( n1852 , n1847 , n1851 ); 
or ( n1853 , n1841 , n1852 ); 
not ( n1854 , n1838 ); 
nand ( n1855 , n388 , n392 ); 
not ( n1856 , n1855 ); 
and ( n1857 , n1854 , n1856 , n1800 ); 
not ( n1858 , n388 ); 
nor ( n1859 , n1858 , n392 ); 
not ( n1860 , n1859 ); 
buf ( n1861 , n1860 ); 
nor ( n1862 , n1835 , n1861 ); 
and ( n1863 , n785 , n1862 ); 
nor ( n1864 , n1857 , n1863 ); 
or ( n1865 , n1864 , n822 ); 
nand ( n1866 , n1853 , n1865 , n1650 ); 
nand ( n1867 , n386 , n1866 ); 
nand ( n1868 , n1844 , n1867 ); 
nand ( n1869 , n1643 , n387 ); 
and ( n1870 , n1869 , n1574 ); 
not ( n1871 , n1669 ); 
nor ( n1872 , n1870 , n1871 ); 
nand ( n1873 , n1524 , n1872 ); 
nand ( n1874 , n1873 , n1589 ); 
not ( n1875 , n1841 ); 
nand ( n1876 , n761 , n1059 ); 
nand ( n1877 , n1875 , n1039 , n1876 , n1744 ); 
not ( n1878 , n1727 ); 
or ( n1879 , n1878 , n1744 ); 
and ( n1880 , n993 , n396 ); 
nand ( n1881 , n1880 , n416 ); 
nand ( n1882 , n1879 , n1881 ); 
nor ( n1883 , n1388 , n794 ); 
nand ( n1884 , n1882 , n1883 ); 
nor ( n1885 , n842 , n1290 , n1330 ); 
or ( n1886 , n1723 , n1885 ); 
nand ( n1887 , n1886 , n396 ); 
nand ( n1888 , n1880 , n1705 ); 
nand ( n1889 , n1887 , n1888 ); 
or ( n1890 , n1289 , n1422 ); 
or ( n1891 , n1425 , n1239 ); 
nand ( n1892 , n1890 , n1891 ); 
nand ( n1893 , n1889 , n1892 , n1214 ); 
nand ( n1894 , n1884 , n1893 ); 
nand ( n1895 , n840 , n402 , n414 ); 
or ( n1896 , n1135 , n913 ); 
nand ( n1897 , n1896 , n995 ); 
and ( n1898 , n777 , n1734 ); 
and ( n1899 , n1895 , n1897 , n1898 ); 
nor ( n1900 , n1899 , n1744 ); 
nor ( n1901 , n1894 , n1900 ); 
not ( n1902 , n1880 ); 
nor ( n1903 , n1902 , n750 , n414 ); 
and ( n1904 , n1903 , n407 ); 
and ( n1905 , n1882 , n407 ); 
and ( n1906 , n1565 , n1035 , n1033 , n1686 ); 
and ( n1907 , n1031 , n1906 , n1069 ); 
nor ( n1908 , n1907 , n1902 ); 
nor ( n1909 , n1904 , n1905 , n1908 ); 
not ( n1910 , n1881 ); 
or ( n1911 , n1903 , n1910 ); 
buf ( n1912 , n1282 ); 
nand ( n1913 , n1911 , n1912 ); 
nand ( n1914 , n1877 , n1901 , n1909 , n1913 ); 
or ( n1915 , n1855 , n390 ); 
or ( n1916 , n785 , n415 ); 
nand ( n1917 , n1916 , n1855 , n416 ); 
nand ( n1918 , n1915 , n1917 ); 
nand ( n1919 , n988 , n1572 ); 
and ( n1920 , n1643 , n1648 ); 
and ( n1921 , n1671 , n1552 ); 
nor ( n1922 , n1920 , n1921 ); 
or ( n1923 , n1919 , n1922 ); 
nor ( n1924 , n1196 , n1496 ); 
and ( n1925 , n1493 , n1924 ); 
nand ( n1926 , n1674 , n1572 ); 
nor ( n1927 , n1926 , n1667 ); 
and ( n1928 , n394 , n1927 ); 
nor ( n1929 , n1925 , n1928 , n1521 ); 
nand ( n1930 , n1923 , n1929 ); 
nor ( n1931 , n1854 , n404 ); 
nand ( n1932 , n1860 , n407 ); 
or ( n1933 , n1931 , n1932 ); 
not ( n1934 , n390 ); 
nand ( n1935 , n1934 , n1859 ); 
nand ( n1936 , n1933 , n1935 ); 
not ( n1937 , n1616 ); 
or ( n1938 , n1937 , n1633 ); 
nand ( n1939 , n1938 , n385 ); 
not ( n1940 , n1922 ); 
and ( n1941 , n1940 , n1673 ); 
nor ( n1942 , n1941 , n1927 ); 
or ( n1943 , n1942 , n394 ); 
not ( n1944 , n1166 ); 
buf ( n1945 , n1496 ); 
or ( n1946 , n1944 , n1945 ); 
nand ( n1947 , n1943 , n1946 ); 
nand ( n1948 , n403 , n901 ); 
or ( n1949 , n1948 , n918 , n1540 ); 
and ( n1950 , n918 , n406 ); 
or ( n1951 , n1197 , n406 ); 
nand ( n1952 , n1951 , n883 ); 
nor ( n1953 , n1950 , n1952 , n1948 ); 
or ( n1954 , n1953 , n775 ); 
nand ( n1955 , n1949 , n1954 ); 
and ( n1956 , n401 , n1952 ); 
not ( n1957 , n883 ); 
not ( n1958 , n44 ); 
and ( n1959 , n1957 , n1958 ); 
nor ( n1960 , n1956 , n1959 ); 
or ( n1961 , n1960 , n1948 ); 
not ( n1962 , n1069 ); 
and ( n1963 , n1898 , n1962 ); 
and ( n1964 , n1948 , n406 ); 
nor ( n1965 , n1963 , n1964 ); 
nand ( n1966 , n1961 , n1965 ); 
nor ( n1967 , n1540 , n1064 ); 
buf ( n1968 , n1967 ); 
and ( n1969 , n394 , n1968 ); 
not ( n1970 , n394 ); 
not ( n1971 , n1609 ); 
and ( n1972 , n1971 , n735 ); 
and ( n1973 , n1970 , n1972 ); 
nor ( n1974 , n1969 , n1973 ); 
nand ( n1975 , n768 , n392 , n1489 ); 
nor ( n1976 , n1974 , n1975 ); 
or ( n1977 , n1976 , n1290 ); 
buf ( n1978 , n1972 ); 
and ( n1979 , n1978 , n759 , n359 ); 
and ( n1980 , n1968 , n344 , n394 ); 
nor ( n1981 , n1979 , n1980 ); 
or ( n1982 , n1975 , n1981 ); 
nor ( n1983 , n1978 , n394 ); 
and ( n1984 , n1967 , n901 ); 
buf ( n1985 , n1984 ); 
nor ( n1986 , n1565 , n1855 , n718 ); 
nand ( n1987 , n1983 , n1985 , n768 , n1986 ); 
nand ( n1988 , n1977 , n1982 , n1987 ); 
not ( n1989 , n822 ); 
nand ( n1990 , n1989 , n1031 ); 
buf ( n1991 , n901 ); 
nand ( n1992 , n1990 , n1991 , n1699 ); 
nand ( n1993 , n1992 , n1565 ); 
nand ( n1994 , n768 , n1489 , n1035 ); 
or ( n1995 , n1981 , n1994 ); 
nor ( n1996 , n1974 , n1994 ); 
or ( n1997 , n1996 , n1330 ); 
nand ( n1998 , n1995 , n1997 ); 
and ( n1999 , n1978 , n759 , n373 ); 
and ( n2000 , n1968 , n44 , n394 ); 
nor ( n2001 , n1999 , n2000 ); 
or ( n2002 , n2001 , n1994 ); 
or ( n2003 , n1996 , n1214 ); 
nand ( n2004 , n2002 , n2003 ); 
not ( n2005 , n1035 ); 
not ( n2006 , n1667 ); 
and ( n2007 , n2005 , n2006 ); 
nor ( n2008 , n2007 , n281 ); 
not ( n2009 , n2008 ); 
not ( n2010 , n392 ); 
not ( n2011 , n1927 ); 
or ( n2012 , n2010 , n2011 ); 
nand ( n2013 , n2012 , n412 ); 
nand ( n2014 , n2009 , n2013 ); 
or ( n2015 , n2001 , n1975 ); 
or ( n2016 , n1976 , n751 ); 
nand ( n2017 , n2015 , n2016 ); 
or ( n2018 , n1155 , n846 ); 
nand ( n2019 , n2018 , n1137 ); 
and ( n2020 , n729 , n2019 ); 
and ( n2021 , n945 , n329 ); 
nor ( n2022 , n2020 , n2021 ); 
or ( n2023 , n2022 , n1945 ); 
or ( n2024 , n729 , n1991 ); 
nand ( n2025 , n2023 , n2024 , n761 ); 
not ( n2026 , n1082 ); 
and ( n2027 , n727 , n1003 ); 
nor ( n2028 , n2027 , n393 ); 
nor ( n2029 , n2026 , n1945 , n2028 ); 
or ( n2030 , n2029 , n846 ); 
and ( n2031 , n1991 , n846 , n1971 ); 
nor ( n2032 , n846 , n857 , n395 ); 
nor ( n2033 , n2031 , n2032 ); 
nand ( n2034 , n2030 , n2033 ); 
nor ( n2035 , n1932 , n404 ); 
not ( n2036 , n2035 ); 
not ( n2037 , n24 ); 
and ( n2038 , n1339 , n2037 , n2 ); 
nor ( n2039 , n2038 , n1912 ); 
or ( n2040 , n2036 , n2039 ); 
not ( n2041 , n417 ); 
and ( n2042 , n2041 , n1114 ); 
and ( n2043 , n409 , n417 ); 
nor ( n2044 , n2042 , n2043 ); 
or ( n2045 , n1256 , n388 ); 
nand ( n2046 , n2045 , n1935 ); 
and ( n2047 , n2046 , n1835 ); 
and ( n2048 , n1856 , n404 ); 
nor ( n2049 , n2047 , n2048 ); 
or ( n2050 , n2044 , n2049 ); 
not ( n2051 , n1861 ); 
or ( n2052 , n1030 , n2051 ); 
nand ( n2053 , n2040 , n2050 , n2052 ); 
or ( n2054 , n388 , n1026 ); 
nand ( n2055 , n2054 , n1915 ); 
and ( n2056 , n2055 , n1801 ); 
and ( n2057 , n2051 , n415 ); 
nor ( n2058 , n2056 , n2057 ); 
or ( n2059 , n2058 , n2044 ); 
or ( n2060 , n1028 , n1856 ); 
not ( n2061 , n1878 ); 
nand ( n2062 , n745 , n751 , n2 , n1703 ); 
not ( n2063 , n2062 ); 
or ( n2064 , n2061 , n2063 ); 
nor ( n2065 , n1856 , n782 , n415 ); 
nand ( n2066 , n2064 , n2065 ); 
nand ( n2067 , n2059 , n2060 , n2066 ); 
not ( n2068 , n760 ); 
not ( n2069 , n2068 ); 
not ( n2070 , n373 ); 
not ( n2071 , n1089 ); 
or ( n2072 , n2070 , n2071 ); 
nand ( n2073 , n2072 , n1312 ); 
not ( n2074 , n2073 ); 
or ( n2075 , n2069 , n2074 ); 
not ( n2076 , n1080 ); 
not ( n2077 , n2076 ); 
not ( n2078 , n846 ); 
and ( n2079 , n2077 , n2078 ); 
not ( n2080 , n880 ); 
and ( n2081 , n1088 , n2080 ); 
nor ( n2082 , n2079 , n2081 ); 
nand ( n2083 , n2075 , n2082 ); 
nor ( n2084 , n1070 , n1945 ); 
not ( n2085 , n1265 ); 
and ( n2086 , n2085 , n398 ); 
and ( n2087 , n775 , n882 ); 
nor ( n2088 , n2087 , n403 ); 
nor ( n2089 , n2086 , n2088 ); 
or ( n2090 , n1945 , n2089 ); 
or ( n2091 , n886 , n1650 ); 
nand ( n2092 , n2090 , n2091 , n1070 ); 
not ( n2093 , n1985 ); 
nor ( n2094 , n2093 , n44 ); 
and ( n2095 , n1876 , n1650 ); 
not ( n2096 , n1985 ); 
not ( n2097 , n1009 ); 
nor ( n2098 , n2096 , n2097 ); 
nor ( n2099 , n2096 , n1197 ); 
nor ( n2100 , n2093 , n1044 ); 
and ( n2101 , n846 , n395 ); 
nand ( n2102 , n393 , n901 ); 
nor ( n2103 , n2101 , n2102 ); 
or ( n2104 , n2103 , n857 ); 
or ( n2105 , n1654 , n1609 ); 
and ( n2106 , n1088 , n846 ); 
nor ( n2107 , n2106 , n2032 ); 
nand ( n2108 , n2104 , n2105 , n2107 ); 
not ( n2109 , n283 ); 
and ( n2110 , n1972 , n901 ); 
not ( n2111 , n2110 ); 
nor ( n2112 , n2109 , n2111 ); 
and ( n2113 , n1985 , n164 ); 
or ( n2114 , n44 , n406 ); 
nand ( n2115 , n2114 , n886 ); 
not ( n2116 , n2115 ); 
not ( n2117 , n903 ); 
or ( n2118 , n2116 , n2117 ); 
nand ( n2119 , n2118 , n398 ); 
and ( n2120 , n1991 , n1065 , n406 ); 
or ( n2121 , n344 , n403 ); 
nand ( n2122 , n2121 , n1958 ); 
and ( n2123 , n775 , n2122 ); 
nor ( n2124 , n2123 , n883 ); 
nor ( n2125 , n2120 , n2124 ); 
nand ( n2126 , n2119 , n2125 ); 
not ( n2127 , n106 ); 
nor ( n2128 , n2127 , n2111 ); 
nor ( n2129 , n2111 , n1155 ); 
not ( n2130 , n313 ); 
nor ( n2131 , n2130 , n2111 ); 
not ( n2132 , n85 ); 
nor ( n2133 , n2132 , n2111 ); 
and ( n2134 , n1985 , n73 ); 
not ( n2135 , n151 ); 
nor ( n2136 , n2135 , n2111 ); 
not ( n2137 , n297 ); 
nor ( n2138 , n2137 , n2111 ); 
not ( n2139 , n266 ); 
nor ( n2140 , n2139 , n2111 ); 
not ( n2141 , n267 ); 
nor ( n2142 , n2141 , n2111 ); 
not ( n2143 , n375 ); 
nor ( n2144 , n2143 , n2111 ); 
and ( n2145 , n1985 , n52 ); 
and ( n2146 , n1985 , n163 ); 
and ( n2147 , n1985 , n95 ); 
and ( n2148 , n1985 , n74 ); 
and ( n2149 , n1985 , n32 ); 
and ( n2150 , n1985 , n190 ); 
and ( n2151 , n1985 , n206 ); 
and ( n2152 , n1313 , n373 ); 
nor ( n2153 , n2152 , n1164 ); 
nor ( n2154 , n2111 , n2153 ); 
and ( n2155 , n1985 , n199 ); 
and ( n2156 , n1985 , n181 ); 
not ( n2157 , n331 ); 
nor ( n2158 , n2157 , n2111 ); 
not ( n2159 , n332 ); 
nor ( n2160 , n2159 , n2111 ); 
and ( n2161 , n1985 , n117 ); 
nor ( n2162 , n2111 , n373 ); 
not ( n2163 , n345 ); 
nor ( n2164 , n2163 , n2111 ); 
not ( n2165 , n346 ); 
nor ( n2166 , n2165 , n2111 ); 
and ( n2167 , n1985 , n141 ); 
not ( n2168 , n312 ); 
nor ( n2169 , n2168 , n2111 ); 
and ( n2170 , n1985 , n162 ); 
and ( n2171 , n1985 , n116 ); 
not ( n2172 , n128 ); 
nor ( n2173 , n2172 , n2111 ); 
not ( n2174 , n330 ); 
nor ( n2175 , n2174 , n2111 ); 
not ( n2176 , n282 ); 
nor ( n2177 , n2176 , n2111 ); 
not ( n2178 , n360 ); 
nor ( n2179 , n2178 , n2111 ); 
not ( n2180 , n374 ); 
nor ( n2181 , n2180 , n2111 ); 
and ( n2182 , n1985 , n11 ); 
and ( n2183 , n1985 , n33 ); 
and ( n2184 , n1985 , n53 ); 
not ( n2185 , n129 ); 
nor ( n2186 , n2185 , n2111 ); 
not ( n2187 , n152 ); 
nor ( n2188 , n2187 , n2111 ); 
not ( n2189 , n86 ); 
nor ( n2190 , n2189 , n2111 ); 
and ( n2191 , n1985 , n140 ); 
not ( n2192 , n361 ); 
nor ( n2193 , n2192 , n2111 ); 
and ( n2194 , n1985 , n118 ); 
and ( n2195 , n1985 , n10 ); 
not ( n2196 , n410 ); 
not ( n2197 , n1926 ); 
or ( n2198 , n2196 , n2197 ); 
or ( n2199 , n1260 , n410 ); 
not ( n2200 , n1848 ); 
nand ( n2201 , n2199 , n2200 ); 
nand ( n2202 , n2198 , n2201 ); 
nand ( n2203 , n2200 , n1260 , n821 ); 
not ( n2204 , n2203 ); 
not ( n2205 , n411 ); 
or ( n2206 , n2204 , n2205 ); 
or ( n2207 , n966 , n2203 ); 
nand ( n2208 , n2206 , n2207 ); 
and ( n2209 , n1985 , n139 ); 
nor ( n2210 , n2111 , n1003 , n1313 ); 
and ( n2211 , n1985 , n94 ); 
not ( n2212 , n296 ); 
nor ( n2213 , n2212 , n2111 ); 
and ( n2214 , n1985 , n96 ); 
not ( n2215 , n408 ); 
or ( n2216 , n2008 , n2215 ); 
nand ( n2217 , n2008 , n1687 ); 
nand ( n2218 , n2216 , n2217 , n1682 ); 
not ( n2219 , n417 ); 
not ( n2220 , n1935 ); 
or ( n2221 , n2219 , n2220 ); 
or ( n2222 , n759 , n1935 ); 
nand ( n2223 , n2221 , n2222 ); 
not ( n2224 , n409 ); 
not ( n2225 , n1915 ); 
or ( n2226 , n2224 , n2225 ); 
or ( n2227 , n759 , n1915 ); 
nand ( n2228 , n2226 , n2227 ); 
not ( n2229 , n2102 ); 
not ( n2230 , n2083 ); 
not ( n2231 , n1650 ); 
or ( n2232 , n2230 , n2231 ); 
or ( n2233 , n2229 , n727 ); 
nand ( n2234 , n2232 , n2233 ); 
not ( n2235 , n1659 ); 
nand ( n2236 , n2235 , n1874 , n1939 ); 
patch p0 (.t_0(t_0), .t_1(t_1), .g1(g343), .g2(g43), .g3(g389), .g4(g387), .g5(g393), .g6(g384), .g7(g390), .g8(g404), .g9(g396), .g10(g400), .g11(g405), .g12(g402), .g13(g397), .g14(g394), .g15(g386), .g16(g399), .g17(g392), .g18(g388), .g19(g372), .g20(g358), .g21(g357), .g22(g280), .g23(g264), .g24(g391), .g25(g371), .g26(g23), .g27(g310), .g28(g63), .g29(g414), .g30(g415), .g31(g403), .g32(g406), .g33(g411), .g34(g409), .g35(g398), .g36(g416), .g37(g401), .g38(g385), .g39(g412), .g40(g408), .g41(g413), .g42(g328));
endmodule 

