module patch (t_0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16);
input g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16;
output t_0;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335;

and ( w1 , g1 , w882 );
nor ( w2 , g2 , g3 );
and ( w3 , w1 , w941 );
nor ( w4 , g5 , g6 );
and ( w5 , w4 , w1135 );
not ( w6 , w5 );
and ( w7 , w6 , g8 );
not ( w8 , w7 );
and ( w9 , g4 , w8 );
and ( w10 , w9 , g8 );
not ( w11 , g9 );
and ( w12 , w11 , g5 );
and ( w13 , w12 , w1236 );
and ( w14 , g9 , g5 );
nor ( w15 , g9 , g5 );
nor ( w16 , w14 , w15 );
not ( w17 , w16 );
and ( w18 , w17 , g6 );
and ( w19 , w18 , w465 );
and ( w20 , w19 , g4 );
nor ( w21 , w13 , w20 );
nor ( w22 , w21 , g10 );
and ( w23 , w882 , g3 );
and ( w24 , g5 , w825 );
and ( w25 , w24 , w1236 );
and ( w26 , g2 , g11 );
and ( w27 , w26 , w1180 );
and ( w28 , g1 , g6 );
not ( w29 , w27 );
and ( w30 , w29 , w28 );
nor ( w31 , w25 , w30 );
nor ( w32 , w31 , w2 );
and ( w33 , w32 , w1105 );
and ( w34 , w33 , g13 );
and ( w35 , w34 , g14 );
and ( w36 , g8 , g7 );
and ( w37 , w36 , g6 );
and ( w38 , w37 , g4 );
and ( w39 , w36 , g5 );
and ( w40 , w39 , w882 );
nor ( w41 , g14 , g12 );
not ( w42 , w41 );
and ( w43 , w42 , g5 );
not ( w44 , w43 );
and ( w45 , w44 , g13 );
nor ( w46 , g12 , g15 );
and ( w47 , w46 , g14 );
and ( w48 , w47 , w1280 );
nor ( w49 , w45 , w48 );
and ( w50 , w41 , g13 );
nor ( w51 , w50 , w48 );
not ( w52 , w51 );
and ( w53 , w52 , g5 );
not ( w54 , w53 );
and ( w55 , w54 , g3 );
nor ( w56 , w55 , w2 );
not ( w57 , w49 );
and ( w58 , w57 , w56 );
and ( w59 , w58 , g11 );
and ( w60 , w59 , w825 );
nor ( w61 , g5 , w26 );
and ( w62 , w61 , w28 );
nor ( w63 , w60 , w62 );
nor ( w64 , g3 , w27 );
and ( w65 , g15 , g14 );
nor ( w66 , w65 , g16 );
not ( w67 , w66 );
and ( w68 , w67 , w28 );
nor ( w69 , w68 , g12 );
not ( w70 , w69 );
and ( w71 , w70 , g6 );
and ( w72 , w71 , w1280 );
nor ( w73 , w64 , w72 );
and ( w74 , w73 , w1105 );
not ( w75 , w74 );
and ( w76 , w75 , w28 );
and ( w77 , w76 , w941 );
not ( w78 , w77 );
and ( w79 , w63 , w78 );
and ( w80 , w79 , w1258 );
nor ( w81 , w80 , w2 );
and ( w82 , w81 , g6 );
nor ( w83 , w40 , w82 );
not ( w84 , w83 );
and ( w85 , w84 , w36 );
and ( w86 , w85 , g4 );
and ( w87 , g4 , g1 );
and ( w88 , w87 , w882 );
and ( w89 , w88 , w941 );
and ( w90 , g1 , w56 );
and ( w91 , w90 , w882 );
and ( w92 , w91 , g7 );
and ( w93 , g5 , w23 );
and ( w94 , g8 , w1135 );
not ( w95 , w93 );
and ( w96 , w95 , w94 );
nor ( w97 , w92 , w96 );
nor ( w98 , w97 , g6 );
and ( w99 , w62 , w941 );
nor ( w100 , w23 , g1 );
and ( w101 , w100 , g11 );
nor ( w102 , w99 , w101 );
not ( w103 , w82 );
and ( w104 , w102 , w103 );
not ( w105 , w104 );
and ( w106 , w105 , g7 );
nor ( w107 , w98 , w106 );
not ( w108 , w107 );
and ( w109 , w108 , g8 );
and ( w110 , w109 , w1258 );
and ( w111 , w110 , w1280 );
and ( w112 , w111 , w1051 );
and ( w113 , w112 , w48 );
nor ( w114 , g8 , g7 );
nor ( w115 , w36 , w114 );
nor ( w116 , w115 , g16 );
and ( w117 , w116 , g1 );
and ( w118 , w117 , g5 );
and ( w119 , w118 , w882 );
and ( w120 , w119 , w941 );
and ( w121 , w120 , w1236 );
nor ( w122 , g13 , w23 );
and ( w123 , w122 , g7 );
and ( w124 , w123 , w1236 );
not ( w125 , w26 );
and ( w126 , w125 , w28 );
and ( w127 , w126 , w941 );
nor ( w128 , w127 , w101 );
nor ( w129 , w128 , g13 );
and ( w130 , w129 , w1135 );
and ( w131 , w130 , w1180 );
nor ( w132 , w124 , w131 );
and ( w133 , g1 , g5 );
and ( w134 , w133 , w882 );
and ( w135 , w134 , w1280 );
and ( w136 , w135 , w1135 );
and ( w137 , w136 , w1236 );
and ( w138 , w62 , w1135 );
nor ( w139 , w137 , w138 );
nor ( w140 , w139 , w2 );
and ( w141 , g5 , g3 );
not ( w142 , w141 );
and ( w143 , w142 , g7 );
and ( w144 , w143 , w1236 );
and ( w145 , w1180 , g3 );
not ( w146 , w145 );
and ( w147 , w146 , g11 );
and ( w148 , w147 , w825 );
and ( w149 , w148 , w1135 );
and ( w150 , w149 , w941 );
nor ( w151 , w144 , w150 );
nor ( w152 , w151 , g13 );
and ( w153 , w152 , w669 );
nor ( w154 , w140 , w153 );
nor ( w155 , w154 , g12 );
and ( w156 , w155 , w1051 );
and ( w157 , w156 , w1280 );
and ( w158 , w157 , w669 );
and ( w159 , w158 , w1258 );
and ( w160 , w159 , g14 );
not ( w161 , w160 );
and ( w162 , w132 , w161 );
not ( w163 , w162 );
and ( w164 , w163 , g4 );
and ( w165 , w164 , w1051 );
nor ( w166 , g13 , g5 );
and ( w167 , w166 , g7 );
and ( w168 , g5 , w1280 );
and ( w169 , w168 , w825 );
and ( w170 , w169 , w1236 );
nor ( w171 , w170 , w28 );
nor ( w172 , w171 , g7 );
and ( w173 , w172 , w1280 );
and ( w174 , w173 , w941 );
and ( w175 , w2 , g1 );
nor ( w176 , w175 , w174 );
not ( w177 , w176 );
and ( w178 , w177 , g5 );
and ( w179 , w178 , w1280 );
and ( w180 , w179 , w1135 );
nor ( w181 , w174 , w180 );
nor ( w182 , w181 , g6 );
nor ( w183 , g5 , w173 );
nor ( w184 , w183 , g7 );
and ( w185 , w184 , w1280 );
and ( w186 , w185 , g6 );
nor ( w187 , w182 , w186 );
not ( w188 , w167 );
and ( w189 , w188 , w187 );
nor ( w190 , w189 , g6 );
nor ( w191 , w190 , w186 );
and ( w192 , w194 , g4 );
and ( w193 , w192 , w465 );
not ( w194 , w191 );
and ( w195 , w194 , g10 );
and ( w196 , w195 , g4 );
and ( w197 , w196 , w669 );
and ( w198 , w197 , w1258 );
and ( w199 , w198 , g14 );
nor ( w200 , w193 , w199 );
nor ( w201 , w200 , g8 );
and ( w202 , w201 , w1258 );
and ( w203 , w202 , g14 );
and ( w204 , g15 , w203 );
nor ( w205 , w165 , w204 );
nor ( w206 , w205 , g8 );
and ( w207 , w206 , g14 );
nor ( w208 , w207 , g7 );
not ( w209 , w208 );
and ( w210 , w209 , g8 );
and ( w211 , w210 , g13 );
nor ( w212 , w207 , w211 );
and ( w213 , w212 , w314 );
nor ( w214 , w213 , w104 );
and ( w215 , w214 , w1105 );
and ( w216 , w215 , g13 );
and ( w217 , w216 , w1282 );
nor ( w218 , g13 , g8 );
and ( w219 , w218 , g7 );
nor ( w220 , w219 , w94 );
nor ( w221 , w220 , g1 );
and ( w222 , w221 , w1180 );
and ( w223 , w222 , w1236 );
and ( w224 , w223 , g4 );
not ( w225 , w4 );
and ( w226 , w225 , g4 );
and ( w227 , w36 , w1280 );
and ( w228 , w227 , g5 );
and ( w229 , w228 , w1236 );
and ( w230 , w227 , g6 );
and ( w231 , w1280 , g7 );
nor ( w232 , w231 , w5 );
not ( w233 , w232 );
and ( w234 , w233 , g8 );
not ( w235 , w234 );
and ( w236 , w235 , g14 );
nor ( w237 , w236 , g13 );
and ( w238 , w237 , g15 );
and ( w239 , w238 , g14 );
nor ( w240 , w207 , w36 );
not ( w241 , w240 );
and ( w242 , w241 , g16 );
not ( w243 , w212 );
and ( w244 , w243 , g12 );
nor ( w245 , w242 , w244 );
and ( w246 , w285 , w245 );
nor ( w247 , w114 , w7 );
nor ( w248 , w247 , g5 );
nor ( w249 , w248 , g16 );
and ( w250 , w249 , w825 );
nor ( w251 , w250 , g6 );
and ( w252 , w825 , g6 );
nor ( w253 , w251 , w252 );
and ( w254 , w28 , g7 );
and ( w255 , w254 , g8 );
nor ( w256 , w114 , w255 );
nor ( w257 , w256 , w252 );
not ( w258 , w257 );
and ( w259 , w258 , g6 );
not ( w260 , w259 );
and ( w261 , w260 , g12 );
and ( w262 , w253 , w261 );
and ( w263 , w262 , w669 );
and ( w264 , w263 , w1135 );
and ( w265 , g8 , w253 );
and ( w266 , w265 , g7 );
nor ( w267 , w264 , w266 );
and ( w268 , w253 , w1180 );
and ( w269 , w268 , w566 );
and ( w270 , w269 , w1236 );
and ( w271 , w270 , w941 );
not ( w272 , w271 );
and ( w273 , w267 , w272 );
nor ( w274 , w273 , w2 );
and ( w275 , w274 , g12 );
and ( w276 , w275 , g10 );
and ( w277 , w276 , g4 );
and ( w278 , w431 , w256 );
not ( w279 , w278 );
and ( w280 , w279 , g12 );
nor ( w281 , w280 , w207 );
and ( w282 , w281 , w314 );
not ( w283 , w242 );
and ( w284 , w283 , w282 );
not ( w285 , w239 );
and ( w286 , w284 , w285 );
and ( w287 , g5 , w566 );
and ( w288 , w287 , w882 );
and ( w289 , w288 , w825 );
and ( w290 , w302 , w71 );
nor ( w291 , w289 , w290 );
not ( w292 , w291 );
and ( w293 , w292 , g15 );
and ( w294 , w293 , g14 );
nor ( w295 , w294 , g16 );
nor ( w296 , w295 , w23 );
nor ( w297 , w296 , w82 );
not ( w298 , w297 );
and ( w299 , w298 , g6 );
and ( w300 , w1280 , w299 );
nor ( w301 , w300 , g12 );
not ( w302 , w288 );
and ( w303 , w302 , w28 );
nor ( w304 , w289 , w303 );
not ( w305 , w304 );
and ( w306 , w305 , g6 );
not ( w307 , w301 );
and ( w308 , w307 , w306 );
and ( w309 , w308 , w961 );
nor ( w310 , w309 , w82 );
nor ( w311 , w286 , w310 );
nor ( w312 , w311 , w207 );
and ( w313 , w246 , w312 );
not ( w314 , w114 );
and ( w315 , w313 , w314 );
nor ( w316 , w315 , w310 );
nor ( w317 , w316 , w207 );
not ( w318 , w317 );
and ( w319 , w230 , w318 );
and ( w320 , w319 , g16 );
nor ( w321 , g1 , w2 );
nor ( w322 , w321 , w175 );
nor ( w323 , w322 , g13 );
and ( w324 , w323 , g5 );
and ( w325 , w324 , g7 );
nor ( w326 , w325 , w5 );
not ( w327 , w326 );
and ( w328 , w327 , g8 );
and ( w329 , w328 , g15 );
and ( w330 , w329 , w1280 );
and ( w331 , w330 , w1258 );
and ( w332 , w331 , w1236 );
not ( w333 , w332 );
and ( w334 , w333 , w317 );
not ( w335 , w334 );
and ( w336 , w335 , g14 );
and ( w337 , w336 , w961 );
nor ( w338 , g16 , g9 );
and ( w339 , w338 , g5 );
and ( w340 , w339 , w1236 );
nor ( w341 , w340 , w306 );
nor ( w342 , w115 , w341 );
and ( w343 , w268 , w1236 );
and ( w344 , w343 , g13 );
nor ( w345 , w344 , w207 );
not ( w346 , w342 );
and ( w347 , w346 , w345 );
and ( w348 , w347 , w465 );
nor ( w349 , w322 , g16 );
and ( w350 , w349 , g5 );
and ( w351 , w350 , w1236 );
nor ( w352 , w351 , w306 );
and ( w353 , w354 , w114 );
not ( w354 , w352 );
and ( w355 , w354 , g7 );
and ( w356 , w355 , g8 );
and ( w357 , g8 , w5 );
nor ( w358 , w357 , w207 );
not ( w359 , w356 );
and ( w360 , w359 , w358 );
and ( w361 , w360 , w345 );
not ( w362 , w361 );
and ( w363 , w362 , g13 );
nor ( w364 , w363 , w207 );
not ( w365 , w353 );
and ( w366 , w365 , w364 );
nor ( w367 , w366 , w23 );
and ( w368 , w367 , g12 );
and ( w369 , w368 , g4 );
and ( w370 , w669 , g7 );
nor ( w371 , w370 , w94 );
nor ( w372 , w371 , g5 );
and ( w373 , w372 , w566 );
and ( w374 , w373 , w825 );
and ( w375 , w374 , w1236 );
and ( w376 , w375 , w1280 );
and ( w377 , w376 , g4 );
and ( w378 , w376 , g10 );
and ( w379 , w378 , g4 );
nor ( w380 , w24 , w82 );
and ( w381 , w458 , g4 );
and ( w382 , w381 , w465 );
and ( w383 , w24 , g10 );
nor ( w384 , w383 , w82 );
not ( w385 , w384 );
and ( w386 , w385 , g4 );
and ( w387 , g4 , w5 );
and ( w388 , w168 , g4 );
and ( w389 , w388 , g7 );
nor ( w390 , w387 , w389 );
nor ( w391 , w390 , g1 );
and ( w392 , w391 , w941 );
and ( w393 , w392 , g8 );
and ( w394 , w393 , g15 );
and ( w395 , w394 , w1280 );
and ( w396 , w395 , w1258 );
and ( w397 , w396 , g14 );
and ( w398 , w262 , g4 );
and ( w399 , w398 , w465 );
nor ( w400 , w399 , w277 );
and ( w401 , w400 , w413 );
not ( w402 , w401 );
and ( w403 , w402 , w114 );
and ( w404 , w271 , g4 );
and ( w405 , w404 , g13 );
nor ( w406 , w405 , w207 );
nor ( w407 , w10 , w207 );
and ( w408 , w406 , w407 );
and ( w409 , w398 , g8 );
and ( w410 , w409 , g7 );
and ( w411 , w410 , w465 );
nor ( w412 , w411 , w277 );
not ( w413 , w207 );
and ( w414 , w412 , w413 );
and ( w415 , w408 , w414 );
nor ( w416 , w415 , g16 );
and ( w417 , w416 , w825 );
and ( w418 , w417 , w465 );
nor ( w419 , w418 , w277 );
nor ( w420 , w419 , w2 );
and ( w421 , w420 , g12 );
and ( w422 , w421 , w1236 );
not ( w423 , w312 );
and ( w424 , g4 , w423 );
and ( w425 , w424 , g14 );
and ( w426 , g4 , w82 );
and ( w427 , w426 , w114 );
and ( w428 , g4 , w255 );
and ( w429 , w428 , g13 );
nor ( w430 , w427 , w429 );
not ( w431 , w277 );
and ( w432 , w430 , w431 );
not ( w433 , w432 );
and ( w434 , w433 , g12 );
nor ( w435 , w434 , w207 );
not ( w436 , w425 );
and ( w437 , w436 , w435 );
not ( w438 , w422 );
and ( w439 , w438 , w437 );
not ( w440 , w403 );
and ( w441 , w440 , w439 );
nor ( w442 , w441 , g1 );
nor ( w443 , w442 , w277 );
nor ( w444 , w443 , w2 );
and ( w445 , w444 , g12 );
and ( w446 , w445 , w1236 );
not ( w447 , w446 );
and ( w448 , w447 , w437 );
not ( w449 , w397 );
and ( w450 , w449 , w448 );
nor ( w451 , w450 , g6 );
not ( w452 , w451 );
and ( w453 , w452 , w437 );
not ( w454 , w386 );
and ( w455 , w454 , w453 );
nor ( w456 , w455 , g13 );
and ( w457 , w456 , w114 );
not ( w458 , w380 );
and ( w459 , w458 , w36 );
and ( w460 , w459 , w1280 );
and ( w461 , w460 , g4 );
nor ( w462 , w461 , w207 );
not ( w463 , w462 );
and ( w464 , w463 , g10 );
not ( w465 , g10 );
and ( w466 , w461 , w465 );
nor ( w467 , w464 , w466 );
not ( w468 , w467 );
and ( w469 , w468 , g7 );
and ( w470 , w469 , g16 );
nor ( w471 , w470 , w207 );
not ( w472 , w457 );
and ( w473 , w472 , w471 );
not ( w474 , w473 );
and ( w475 , w474 , g16 );
not ( w476 , w475 );
and ( w477 , w476 , w453 );
not ( w478 , w382 );
and ( w479 , w478 , w477 );
nor ( w480 , w479 , g13 );
and ( w481 , w480 , w114 );
not ( w482 , w481 );
and ( w483 , w482 , w471 );
not ( w484 , w483 );
and ( w485 , w484 , g16 );
not ( w486 , w485 );
and ( w487 , w486 , w453 );
not ( w488 , w379 );
and ( w489 , w488 , w487 );
not ( w490 , w489 );
and ( w491 , w490 , g16 );
not ( w492 , w491 );
and ( w493 , w492 , w453 );
not ( w494 , w377 );
and ( w495 , w494 , w493 );
nor ( w496 , w495 , g10 );
not ( w497 , w496 );
and ( w498 , w497 , w493 );
not ( w499 , w498 );
and ( w500 , w499 , g16 );
not ( w501 , w500 );
and ( w502 , w501 , w453 );
not ( w503 , w369 );
and ( w504 , w503 , w502 );
nor ( w505 , w348 , w504 );
and ( w506 , w505 , w961 );
and ( w507 , w506 , g12 );
not ( w508 , w507 );
and ( w509 , w508 , w502 );
not ( w510 , w337 );
and ( w511 , w510 , w509 );
not ( w512 , w511 );
and ( w513 , w512 , g4 );
nor ( w514 , w320 , w513 );
not ( w515 , w229 );
and ( w516 , w515 , w514 );
not ( w517 , w516 );
and ( w518 , w517 , g4 );
and ( w519 , w518 , g7 );
and ( w520 , w519 , w1105 );
and ( w521 , w520 , w961 );
and ( w522 , w521 , g16 );
nor ( w523 , w522 , w513 );
not ( w524 , w226 );
and ( w525 , w524 , w523 );
nor ( w526 , w525 , g13 );
and ( w527 , w526 , w114 );
not ( w528 , w527 );
and ( w529 , w528 , w523 );
nor ( w530 , w529 , g12 );
and ( w531 , w530 , w961 );
and ( w532 , w531 , g16 );
nor ( w533 , w532 , w513 );
not ( w534 , w224 );
and ( w535 , w534 , w533 );
nor ( w536 , w535 , w23 );
and ( w537 , w536 , g16 );
nor ( w538 , w537 , w513 );
not ( w539 , w217 );
and ( w540 , w539 , w538 );
not ( w541 , w121 );
and ( w542 , w541 , w540 );
nor ( w543 , w93 , w371 );
and ( w544 , w543 , w1236 );
not ( w545 , w544 );
and ( w546 , w545 , w540 );
nor ( w547 , w546 , g12 );
and ( w548 , w547 , g13 );
and ( w549 , w548 , w1282 );
not ( w550 , w549 );
and ( w551 , w550 , w538 );
and ( w552 , w542 , w551 );
nor ( w553 , w552 , g12 );
and ( w554 , w553 , g13 );
and ( w555 , w554 , w1282 );
not ( w556 , w555 );
and ( w557 , w556 , w538 );
not ( w558 , w113 );
and ( w559 , w558 , w557 );
not ( w560 , w559 );
and ( w561 , w560 , g4 );
nor ( w562 , w89 , w561 );
not ( w563 , w562 );
and ( w564 , w563 , w114 );
nor ( w565 , w23 , g5 );
not ( w566 , g3 );
and ( w567 , w566 , g1 );
nor ( w568 , g1 , g5 );
nor ( w569 , w567 , w568 );
nor ( w570 , w569 , w2 );
nor ( w571 , w565 , w570 );
nor ( w572 , w571 , w371 );
and ( w573 , w572 , g4 );
nor ( w574 , w573 , w207 );
nor ( w575 , w574 , g6 );
nor ( w576 , w575 , w561 );
not ( w577 , w576 );
and ( w578 , w577 , g16 );
nor ( w579 , w578 , w561 );
not ( w580 , w564 );
and ( w581 , w580 , w579 );
nor ( w582 , w581 , g6 );
nor ( w583 , w582 , w561 );
not ( w584 , w583 );
and ( w585 , w584 , g16 );
nor ( w586 , w585 , w561 );
not ( w587 , w86 );
and ( w588 , w587 , w586 );
nor ( w589 , w588 , w2 );
and ( w590 , w589 , g7 );
not ( w591 , w590 );
and ( w592 , w591 , w586 );
not ( w593 , w592 );
and ( w594 , w593 , g16 );
nor ( w595 , w594 , w561 );
not ( w596 , w38 );
and ( w597 , w596 , w595 );
not ( w598 , w597 );
and ( w599 , w598 , g16 );
nor ( w600 , w599 , w561 );
not ( w601 , w35 );
and ( w602 , w601 , w600 );
and ( w603 , w23 , w602 );
not ( w604 , w603 );
and ( w605 , w604 , g9 );
and ( w606 , w605 , g10 );
and ( w607 , w606 , w1105 );
and ( w608 , w607 , g13 );
and ( w609 , w608 , g14 );
not ( w610 , w609 );
and ( w611 , w610 , w600 );
not ( w612 , w611 );
and ( w613 , w612 , g5 );
nor ( w614 , w613 , g6 );
and ( w615 , g9 , g10 );
not ( w616 , w614 );
and ( w617 , w616 , w615 );
and ( w618 , w617 , g4 );
and ( w619 , w1180 , g7 );
nor ( w620 , g9 , g10 );
nor ( w621 , w620 , w615 );
and ( w622 , w1144 , g1 );
and ( w623 , w622 , g5 );
and ( w624 , w623 , w882 );
and ( w625 , w624 , w941 );
and ( w626 , w625 , w114 );
nor ( w627 , w619 , w626 );
not ( w628 , w627 );
and ( w629 , w628 , g4 );
and ( w630 , w1144 , g4 );
and ( w631 , w565 , g4 );
not ( w632 , w631 );
and ( w633 , w632 , w600 );
nor ( w634 , w633 , g6 );
not ( w635 , w620 );
and ( w636 , w635 , w611 );
not ( w637 , w636 );
and ( w638 , w637 , g5 );
and ( w639 , w638 , w1236 );
and ( w640 , g9 , w1180 );
not ( w641 , w640 );
and ( w642 , w641 , w306 );
and ( w643 , w642 , w961 );
and ( w644 , w30 , w941 );
nor ( w645 , w643 , w644 );
nor ( w646 , w645 , g10 );
nor ( w647 , w646 , w615 );
not ( w648 , w647 );
and ( w649 , w648 , g6 );
nor ( w650 , w639 , w649 );
not ( w651 , w650 );
and ( w652 , w651 , g4 );
not ( w653 , w652 );
and ( w654 , w653 , w600 );
not ( w655 , w654 );
and ( w656 , w655 , w114 );
and ( w657 , w656 , w1105 );
and ( w658 , w657 , w1258 );
and ( w659 , w658 , g13 );
and ( w660 , w659 , g14 );
not ( w661 , w660 );
and ( w662 , w661 , w600 );
not ( w663 , w634 );
and ( w664 , w663 , w662 );
not ( w665 , w664 );
and ( w666 , w665 , g7 );
not ( w667 , w666 );
and ( w668 , w667 , w662 );
not ( w669 , g8 );
and ( w670 , w669 , g13 );
and ( w671 , w670 , g14 );
not ( w672 , w668 );
and ( w673 , w672 , w671 );
not ( w674 , w673 );
and ( w675 , w674 , w600 );
not ( w676 , w630 );
and ( w677 , w676 , w675 );
nor ( w678 , w677 , g5 );
not ( w679 , w150 );
and ( w680 , w679 , w600 );
not ( w681 , w680 );
and ( w682 , w681 , g11 );
nor ( w683 , w682 , w62 );
not ( w684 , w683 );
and ( w685 , w684 , g4 );
not ( w686 , w685 );
and ( w687 , w686 , w675 );
nor ( w688 , w687 , w2 );
and ( w689 , w688 , g6 );
not ( w690 , w689 );
and ( w691 , w690 , w675 );
nor ( w692 , w691 , g8 );
and ( w693 , w692 , w1105 );
and ( w694 , w693 , g13 );
and ( w695 , w694 , g14 );
not ( w696 , w695 );
and ( w697 , w696 , w600 );
not ( w698 , w678 );
and ( w699 , w698 , w697 );
not ( w700 , w699 );
and ( w701 , w700 , w114 );
and ( w702 , w701 , g6 );
not ( w703 , w702 );
and ( w704 , w703 , w675 );
not ( w705 , w704 );
and ( w706 , w705 , g13 );
and ( w707 , w706 , g14 );
not ( w708 , w707 );
and ( w709 , w708 , w600 );
not ( w710 , w629 );
and ( w711 , w710 , w709 );
nor ( w712 , w711 , g6 );
not ( w713 , w712 );
and ( w714 , w713 , w709 );
not ( w715 , w714 );
and ( w716 , w715 , w671 );
not ( w717 , w716 );
and ( w718 , w717 , w600 );
not ( w719 , w618 );
and ( w720 , w719 , w718 );
not ( w721 , w720 );
and ( w722 , w721 , g7 );
and ( w723 , w722 , g8 );
not ( w724 , w723 );
and ( w725 , w724 , w718 );
not ( w726 , w725 );
and ( w727 , w726 , g13 );
and ( w728 , w727 , g14 );
not ( w729 , w728 );
and ( w730 , w729 , w600 );
and ( w731 , w763 , w730 );
and ( w732 , w731 , w1236 );
not ( w733 , w732 );
and ( w734 , w733 , w615 );
and ( w735 , w734 , g4 );
not ( w736 , w735 );
and ( w737 , w736 , w718 );
not ( w738 , w737 );
and ( w739 , w738 , g7 );
and ( w740 , w739 , g8 );
not ( w741 , w740 );
and ( w742 , w741 , w718 );
not ( w743 , w742 );
and ( w744 , w743 , g13 );
and ( w745 , w744 , g14 );
not ( w746 , w745 );
and ( w747 , w746 , w600 );
not ( w748 , w22 );
and ( w749 , w748 , w747 );
not ( w750 , w749 );
and ( w751 , w750 , g4 );
and ( w752 , w751 , g7 );
and ( w753 , w752 , g8 );
not ( w754 , w753 );
and ( w755 , w754 , w718 );
not ( w756 , w10 );
and ( w757 , w756 , w755 );
not ( w758 , w757 );
and ( w759 , w758 , g13 );
and ( w760 , w759 , g14 );
not ( w761 , w760 );
and ( w762 , w761 , w600 );
not ( w763 , w3 );
and ( w764 , w763 , w762 );
nor ( w765 , g1 , w371 );
not ( w766 , w765 );
and ( w767 , w766 , w762 );
not ( w768 , g11 );
and ( w769 , w767 , w768 );
nor ( w770 , g5 , g3 );
and ( w771 , w770 , w941 );
not ( w772 , w771 );
and ( w773 , w23 , w772 );
nor ( w774 , w773 , w371 );
and ( w775 , w774 , w1180 );
not ( w776 , w775 );
and ( w777 , w776 , w762 );
not ( w778 , w777 );
and ( w779 , w778 , g1 );
not ( w780 , w779 );
and ( w781 , w780 , w762 );
not ( w782 , w781 );
and ( w783 , w782 , g11 );
not ( w784 , w783 );
and ( w785 , w784 , w762 );
and ( w786 , w785 , g6 );
nor ( w787 , w769 , w786 );
and ( w788 , w787 , g4 );
and ( w789 , w788 , w1105 );
not ( w790 , w789 );
and ( w791 , w790 , w762 );
and ( w792 , w762 , w1040 );
and ( w793 , w792 , g2 );
nor ( w794 , w793 , w371 );
nor ( w795 , w794 , g6 );
and ( w796 , w61 , w825 );
and ( w797 , w941 , w796 );
nor ( w798 , w175 , w797 );
nor ( w799 , w798 , w371 );
not ( w800 , w799 );
and ( w801 , w800 , w762 );
and ( w802 , w801 , g6 );
nor ( w803 , w795 , w802 );
and ( w804 , w803 , w1180 );
not ( w805 , w804 );
and ( w806 , w805 , w762 );
not ( w807 , w806 );
and ( w808 , w807 , g4 );
and ( w809 , w808 , w1105 );
not ( w810 , w809 );
and ( w811 , w810 , w762 );
not ( w812 , w568 );
and ( w813 , w812 , w762 );
and ( w814 , w873 , g4 );
not ( w815 , w371 );
and ( w816 , w814 , w815 );
not ( w817 , w816 );
and ( w818 , w817 , w762 );
not ( w819 , w818 );
and ( w820 , w819 , g6 );
not ( w821 , w820 );
and ( w822 , w821 , w762 );
nor ( w823 , w371 , g3 );
and ( w824 , w823 , g5 );
not ( w825 , g1 );
and ( w826 , w824 , w825 );
and ( w827 , w826 , w882 );
not ( w828 , w827 );
and ( w829 , w828 , w762 );
and ( w830 , w762 , g10 );
and ( w831 , w830 , w1040 );
and ( w832 , w831 , g7 );
nor ( w833 , w288 , w371 );
not ( w834 , w832 );
and ( w835 , w834 , w833 );
and ( w836 , w835 , g1 );
not ( w837 , w836 );
and ( w838 , w837 , w762 );
and ( w839 , w829 , w838 );
not ( w840 , w839 );
and ( w841 , w840 , g12 );
not ( w842 , w841 );
and ( w843 , w842 , w762 );
and ( w844 , g1 , g11 );
nor ( w845 , w220 , g13 );
and ( w846 , w844 , w845 );
not ( w847 , w133 );
and ( w848 , w847 , w845 );
not ( w849 , w848 );
and ( w850 , w849 , w762 );
nor ( w851 , w850 , g6 );
not ( w852 , w851 );
and ( w853 , w852 , w762 );
nor ( w854 , w853 , g13 );
and ( w855 , w854 , g14 );
not ( w856 , w855 );
and ( w857 , w856 , w762 );
not ( w858 , w846 );
and ( w859 , w858 , w857 );
nor ( w860 , w859 , g5 );
and ( w861 , w860 , w1051 );
not ( w862 , w861 );
and ( w863 , w862 , w762 );
not ( w864 , w798 );
and ( w865 , w864 , g6 );
not ( w866 , w865 );
and ( w867 , w866 , w857 );
not ( w868 , w867 );
and ( w869 , w868 , w845 );
not ( w870 , w869 );
and ( w871 , w870 , w762 );
nor ( w872 , w871 , g15 );
not ( w873 , w813 );
and ( w874 , w873 , w845 );
not ( w875 , w874 );
and ( w876 , w875 , w762 );
not ( w877 , w876 );
and ( w878 , w877 , g6 );
not ( w879 , w878 );
and ( w880 , w879 , w762 );
nor ( w881 , g3 , g1 );
not ( w882 , g2 );
and ( w883 , w881 , w882 );
and ( w884 , w926 , g1 );
and ( w885 , w884 , w1236 );
not ( w886 , w885 );
and ( w887 , w886 , w762 );
nor ( w888 , w887 , g13 );
and ( w889 , w941 , w888 );
nor ( w890 , w883 , w889 );
and ( w891 , w890 , g5 );
not ( w892 , w891 );
and ( w893 , w892 , w845 );
not ( w894 , w893 );
and ( w895 , w894 , w762 );
nor ( w896 , w895 , g6 );
not ( w897 , w896 );
and ( w898 , w897 , w762 );
nor ( w899 , w898 , g13 );
not ( w900 , w899 );
and ( w901 , w880 , w900 );
not ( w902 , w901 );
and ( w903 , w902 , g15 );
and ( w904 , w903 , g14 );
not ( w905 , w904 );
and ( w906 , w905 , w762 );
nor ( w907 , w906 , w23 );
and ( w908 , w567 , w771 );
and ( w909 , w908 , g11 );
nor ( w910 , w909 , w796 );
not ( w911 , w910 );
and ( w912 , w911 , w845 );
not ( w913 , w912 );
and ( w914 , w913 , w762 );
not ( w915 , w914 );
and ( w916 , w915 , g6 );
not ( w917 , w916 );
and ( w918 , w917 , w762 );
and ( w919 , w918 , w857 );
nor ( w920 , w919 , g12 );
and ( w921 , w920 , w1051 );
not ( w922 , w921 );
and ( w923 , w922 , w762 );
nor ( w924 , g11 , g3 );
and ( w925 , w924 , g4 );
not ( w926 , w220 );
and ( w927 , w926 , w925 );
not ( w928 , w927 );
and ( w929 , w928 , w762 );
nor ( w930 , w929 , g1 );
not ( w931 , w930 );
and ( w932 , w931 , w762 );
not ( w933 , w932 );
and ( w934 , w933 , g6 );
not ( w935 , w934 );
and ( w936 , w935 , w762 );
not ( w937 , w888 );
and ( w938 , w936 , w937 );
not ( w939 , w938 );
and ( w940 , w939 , g15 );
not ( w941 , w2 );
and ( w942 , w940 , w941 );
and ( w943 , w942 , g4 );
and ( w944 , w943 , g14 );
not ( w945 , w944 );
and ( w946 , w945 , w762 );
nor ( w947 , w946 , g13 );
not ( w948 , w947 );
and ( w949 , w923 , w948 );
nor ( w950 , w949 , w2 );
and ( w951 , w950 , w1280 );
and ( w952 , w951 , g4 );
not ( w953 , w952 );
and ( w954 , w953 , w762 );
not ( w955 , w954 );
and ( w956 , w955 , g14 );
not ( w957 , w956 );
and ( w958 , w957 , w762 );
nor ( w959 , w792 , w371 );
and ( w960 , w959 , w1236 );
not ( w961 , w23 );
and ( w962 , w568 , w961 );
nor ( w963 , w962 , w925 );
not ( w964 , w963 );
and ( w965 , w964 , g4 );
not ( w966 , w965 );
and ( w967 , w571 , w966 );
not ( w968 , w967 );
and ( w969 , w968 , g4 );
not ( w970 , w969 );
and ( w971 , w970 , w762 );
nor ( w972 , w971 , w371 );
and ( w973 , w972 , g6 );
not ( w974 , w973 );
and ( w975 , w974 , w762 );
not ( w976 , w960 );
and ( w977 , w976 , w975 );
nor ( w978 , w977 , g16 );
not ( w979 , w978 );
and ( w980 , w979 , w762 );
nor ( w981 , w980 , g13 );
and ( w982 , w981 , w1282 );
not ( w983 , w982 );
and ( w984 , w983 , w762 );
and ( w985 , w958 , w984 );
not ( w986 , w907 );
and ( w987 , w986 , w985 );
not ( w988 , w987 );
and ( w989 , w988 , g4 );
nor ( w990 , w872 , w989 );
nor ( w991 , w990 , w23 );
not ( w992 , w991 );
and ( w993 , w992 , w985 );
nor ( w994 , w993 , g13 );
and ( w995 , w994 , g4 );
not ( w996 , w995 );
and ( w997 , w996 , w762 );
not ( w998 , w997 );
and ( w999 , w998 , g14 );
not ( w1000 , w999 );
and ( w1001 , w1000 , w762 );
and ( w1002 , w1001 , w984 );
and ( w1003 , w863 , w1002 );
nor ( w1004 , w1003 , w23 );
not ( w1005 , w1004 );
and ( w1006 , w1005 , w985 );
nor ( w1007 , w1006 , g13 );
and ( w1008 , w1007 , g4 );
not ( w1009 , w1008 );
and ( w1010 , w1009 , w762 );
not ( w1011 , w1010 );
and ( w1012 , w1011 , g14 );
not ( w1013 , w1012 );
and ( w1014 , w1013 , w762 );
and ( w1015 , w1014 , w984 );
and ( w1016 , w843 , w1015 );
nor ( w1017 , w792 , w1016 );
and ( w1018 , w1017 , w1236 );
not ( w1019 , w1018 );
and ( w1020 , w1019 , w762 );
and ( w1021 , w1020 , w1015 );
and ( w1022 , w822 , w1021 );
not ( w1023 , w1022 );
and ( w1024 , w1023 , g12 );
not ( w1025 , w1024 );
and ( w1026 , w1025 , w762 );
and ( w1027 , w1026 , w1015 );
and ( w1028 , w811 , w1027 );
nor ( w1029 , w1028 , g14 );
and ( w1030 , w1029 , g13 );
not ( w1031 , w1030 );
and ( w1032 , w1031 , w762 );
and ( w1033 , w1032 , w1015 );
and ( w1034 , w791 , w1033 );
nor ( w1035 , w1034 , g14 );
and ( w1036 , w1035 , g13 );
not ( w1037 , w1036 );
and ( w1038 , w1037 , w762 );
and ( w1039 , w1038 , w1015 );
not ( w1040 , g4 );
and ( w1041 , w1039 , w1040 );
and ( w1042 , w93 , g6 );
and ( w1043 , w1042 , w1280 );
not ( w1044 , w1043 );
and ( w1045 , w1044 , w762 );
not ( w1046 , w1045 );
and ( w1047 , w1046 , w114 );
not ( w1048 , w1047 );
and ( w1049 , w1048 , w762 );
nor ( w1050 , w1049 , g12 );
not ( w1051 , g15 );
and ( w1052 , w1050 , w1051 );
not ( w1053 , w1052 );
and ( w1054 , w1053 , w1039 );
nor ( w1055 , w1054 , g13 );
not ( w1056 , w1055 );
and ( w1057 , w1056 , w762 );
not ( w1058 , w1057 );
and ( w1059 , w1058 , g14 );
not ( w1060 , w1059 );
and ( w1061 , w1060 , w762 );
not ( w1062 , w1042 );
and ( w1063 , w1062 , w762 );
not ( w1064 , w1063 );
and ( w1065 , w1064 , w114 );
not ( w1066 , w1065 );
and ( w1067 , w1066 , w762 );
not ( w1068 , w1067 );
and ( w1069 , w1068 , g13 );
not ( w1070 , w1069 );
and ( w1071 , w1070 , w762 );
and ( w1072 , g5 , g6 );
not ( w1073 , w1072 );
and ( w1074 , w1073 , w762 );
nor ( w1075 , w1074 , g16 );
not ( w1076 , w1075 );
and ( w1077 , w1076 , w762 );
not ( w1078 , w1077 );
and ( w1079 , w1078 , w114 );
not ( w1080 , w1079 );
and ( w1081 , w1080 , w762 );
nor ( w1082 , w1081 , g13 );
not ( w1083 , w1082 );
and ( w1084 , w1083 , w762 );
nor ( w1085 , w1084 , g14 );
not ( w1086 , w1085 );
and ( w1087 , w1071 , w1086 );
nor ( w1088 , w1087 , g12 );
and ( w1089 , w1088 , w1282 );
not ( w1090 , w1089 );
and ( w1091 , w1090 , w1039 );
nor ( w1092 , w1074 , g12 );
and ( w1093 , w1092 , g13 );
and ( w1094 , w1093 , g14 );
not ( w1095 , w1094 );
and ( w1096 , w1095 , w762 );
and ( w1097 , g15 , g6 );
and ( w1098 , w1097 , g5 );
not ( w1099 , w1098 );
and ( w1100 , w1099 , w762 );
nor ( w1101 , w1100 , g13 );
and ( w1102 , w1101 , g14 );
not ( w1103 , w1102 );
and ( w1104 , w1103 , w762 );
not ( w1105 , g12 );
and ( w1106 , w1072 , w1105 );
and ( w1107 , w1106 , w1280 );
not ( w1108 , w1107 );
and ( w1109 , w1108 , w762 );
nor ( w1110 , w1109 , g14 );
and ( w1111 , w1110 , g4 );
not ( w1112 , w1111 );
and ( w1113 , w1112 , w762 );
and ( w1114 , g5 , g12 );
and ( w1115 , g6 , w1114 );
not ( w1116 , w1115 );
and ( w1117 , w1116 , w762 );
not ( w1118 , w1117 );
and ( w1119 , w1118 , g4 );
and ( w1120 , w1119 , w1282 );
not ( w1121 , w1120 );
and ( w1122 , w1113 , w1121 );
nor ( w1123 , w1122 , g14 );
not ( w1124 , w1123 );
and ( w1125 , w1104 , w1124 );
and ( w1126 , w1096 , w1125 );
not ( w1127 , w1126 );
and ( w1128 , w1127 , w114 );
and ( w1129 , w621 , g4 );
not ( w1130 , w1129 );
and ( w1131 , w1130 , w762 );
and ( w1132 , w1131 , g5 );
not ( w1133 , w1132 );
and ( w1134 , w1133 , g8 );
not ( w1135 , g7 );
and ( w1136 , w1134 , w1135 );
not ( w1137 , w1136 );
and ( w1138 , w1137 , w762 );
not ( w1139 , w1138 );
and ( w1140 , w1139 , g13 );
and ( w1141 , w1140 , w94 );
not ( w1142 , w1141 );
and ( w1143 , w1142 , w762 );
not ( w1144 , w621 );
and ( w1145 , w1144 , g5 );
not ( w1146 , w1145 );
and ( w1147 , w1146 , g4 );
not ( w1148 , w1147 );
and ( w1149 , w1148 , w762 );
and ( w1150 , w1149 , w1236 );
not ( w1151 , w1150 );
and ( w1152 , g7 , w1151 );
not ( w1153 , w1152 );
and ( w1154 , w1153 , w762 );
not ( w1155 , w1154 );
and ( w1156 , w1155 , g13 );
and ( w1157 , w1156 , w671 );
not ( w1158 , w1157 );
and ( w1159 , w1158 , w1033 );
and ( w1160 , w1159 , w1236 );
and ( w1161 , w621 , w1180 );
and ( w1162 , w1161 , g4 );
nor ( w1163 , g14 , g13 );
not ( w1164 , w1163 );
and ( w1165 , w1164 , w762 );
not ( w1166 , w925 );
and ( w1167 , w1166 , w762 );
and ( w1168 , w1167 , g6 );
and ( w1169 , w1168 , g5 );
and ( w1170 , w1171 , w94 );
not ( w1171 , w1169 );
and ( w1172 , w1171 , g7 );
and ( w1173 , w1172 , w671 );
not ( w1174 , w1173 );
and ( w1175 , w1174 , w762 );
not ( w1176 , w1170 );
and ( w1177 , w1176 , w1175 );
not ( w1178 , w1177 );
and ( w1179 , w621 , w1178 );
not ( w1180 , g5 );
and ( w1181 , w1179 , w1180 );
and ( w1182 , w1181 , g4 );
not ( w1183 , w1182 );
and ( w1184 , w1183 , w762 );
nor ( w1185 , w1184 , g16 );
not ( w1186 , w1185 );
and ( w1187 , w1186 , w762 );
not ( w1188 , w1187 );
and ( w1189 , w1188 , g13 );
and ( w1190 , w1189 , g14 );
not ( w1191 , w1190 );
and ( w1192 , w1191 , w762 );
and ( w1193 , w1192 , w1039 );
and ( w1194 , w1193 , g6 );
and ( w1195 , w1165 , w1194 );
not ( w1196 , w1162 );
and ( w1197 , w1196 , w1195 );
nor ( w1198 , w1197 , g7 );
and ( w1199 , w1198 , g8 );
and ( w1200 , w1199 , g13 );
not ( w1201 , w1200 );
and ( w1202 , w1201 , w762 );
not ( w1203 , w1195 );
and ( w1204 , w1203 , g4 );
and ( w1205 , w1204 , g7 );
not ( w1206 , w1205 );
and ( w1207 , w1206 , w762 );
not ( w1208 , w1207 );
and ( w1209 , w1208 , g13 );
not ( w1210 , w1209 );
and ( w1211 , w1210 , w1033 );
not ( w1212 , w1211 );
and ( w1213 , w1212 , g14 );
not ( w1214 , w1213 );
and ( w1215 , w1214 , w762 );
and ( w1216 , w1215 , w1033 );
and ( w1217 , w1216 , g6 );
and ( w1218 , w1202 , w1217 );
nor ( w1219 , w1218 , g16 );
not ( w1220 , w1219 );
and ( w1221 , w1220 , w762 );
not ( w1222 , w1221 );
and ( w1223 , w1222 , g14 );
not ( w1224 , w1223 );
and ( w1225 , w1224 , w762 );
and ( w1226 , w1225 , w1033 );
and ( w1227 , w1226 , g6 );
nor ( w1228 , w1160 , w1227 );
not ( w1229 , w1228 );
and ( w1230 , w1143 , w1229 );
not ( w1231 , w1230 );
and ( w1232 , w1231 , g14 );
not ( w1233 , w1232 );
and ( w1234 , w1233 , w762 );
and ( w1235 , w1234 , w1033 );
not ( w1236 , g6 );
and ( w1237 , w1235 , w1236 );
nor ( w1238 , w1237 , w1227 );
nor ( w1239 , w1128 , w1238 );
and ( w1240 , w1091 , w1239 );
and ( w1241 , w1061 , w1240 );
nor ( w1242 , w1041 , w1241 );
not ( w1243 , w1114 );
and ( w1244 , w764 , w1243 );
not ( w1245 , w1244 );
and ( w1246 , w1245 , g6 );
not ( w1247 , w1246 );
and ( w1248 , w1247 , w762 );
nor ( w1249 , g7 , w1242 );
nor ( w1250 , w1248 , w1249 );
nor ( w1251 , w1250 , w1242 );
not ( w1252 , w1251 );
and ( w1253 , w1252 , g13 );
nor ( w1254 , g5 , w1110 );
not ( w1255 , w1254 );
and ( w1256 , w1255 , g6 );
and ( w1257 , w1256 , w36 );
not ( w1258 , g16 );
and ( w1259 , w1257 , w1258 );
not ( w1260 , w1259 );
and ( w1261 , w1260 , w762 );
nor ( w1262 , w1261 , g12 );
and ( w1263 , w1262 , w1280 );
nor ( w1264 , w1263 , w1242 );
nor ( w1265 , w1264 , g14 );
nor ( w1266 , w1265 , w1242 );
not ( w1267 , w1253 );
and ( w1268 , w1267 , w1266 );
not ( w1269 , w1268 );
and ( w1270 , w1269 , g4 );
nor ( w1271 , g8 , w1242 );
and ( w1272 , w1270 , w1303 );
and ( w1273 , w1272 , w1282 );
not ( w1274 , w1273 );
and ( w1275 , w1274 , w762 );
and ( w1276 , w1313 , w1275 );
and ( w1277 , w764 , w1276 );
and ( w1278 , w1277 , w1125 );
nor ( w1279 , w1278 , w1249 );
not ( w1280 , g13 );
and ( w1281 , w1279 , w1280 );
not ( w1282 , g14 );
and ( w1283 , w1282 , w1276 );
and ( w1284 , w1281 , w1298 );
and ( w1285 , w1284 , g6 );
not ( w1286 , w1285 );
and ( w1287 , w1286 , w762 );
and ( w1288 , w1287 , w1276 );
not ( w1289 , w1288 );
and ( w1290 , w1289 , g4 );
and ( w1291 , w1290 , w1303 );
nor ( w1292 , w1291 , g5 );
nor ( w1293 , g13 , w1291 );
nor ( w1294 , g12 , w1293 );
not ( w1295 , w1294 );
and ( w1296 , w1295 , w1276 );
nor ( w1297 , w1292 , w1296 );
not ( w1298 , w1283 );
and ( w1299 , w1297 , w1298 );
not ( w1300 , w1249 );
and ( w1301 , w1299 , w1300 );
nor ( w1302 , w1293 , w1283 );
not ( w1303 , w1271 );
and ( w1304 , w1302 , w1303 );
and ( w1305 , w1301 , w1304 );
and ( w1306 , w1305 , g6 );
not ( w1307 , w1306 );
and ( w1308 , w1307 , w1276 );
not ( w1309 , w1308 );
and ( w1310 , w1309 , g4 );
nor ( w1311 , w1310 , w1291 );
and ( w1312 , w1311 , w762 );
not ( w1313 , w1242 );
and ( w1314 , w1312 , w1313 );
and ( w1315 , w1314 , w762 );
and ( w1316 , w1315 , w1276 );
and ( w1317 , w1316 , w1334 );
and ( w1318 , w1317 , w1315 );
and ( w1319 , w1312 , w1334 );
and ( w1320 , w1318 , w1319 );
and ( w1321 , w1320 , w1334 );
and ( w1322 , w1321 , w1276 );
and ( w1323 , w1322 , w1334 );
and ( w1324 , w1323 , w1315 );
and ( w1325 , w1324 , w1320 );
and ( w1326 , w1316 , w1319 );
and ( w1327 , w1325 , w1326 );
and ( w1328 , w1327 , w1315 );
and ( w1329 , w1328 , w1326 );
and ( w1330 , w1329 , w1320 );
and ( w1331 , w1330 , w1323 );
and ( w1332 , w1331 , w1276 );
and ( w1333 , w1332 , w1334 );
not ( w1334 , w1291 );
and ( w1335 , w1327 , w1334 );
and ( t_0 , w1333 , w1335 );

endmodule
