module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 ; 
output g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
n2920 , n2921 , n2922 ; 
wire t_0 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( n158 , g157 ); 
buf ( n159 , g158 ); 
buf ( n160 , g159 ); 
buf ( n161 , g160 ); 
buf ( n162 , g161 ); 
buf ( n163 , g162 ); 
buf ( n164 , g163 ); 
buf ( n165 , g164 ); 
buf ( n166 , g165 ); 
buf ( n167 , g166 ); 
buf ( n168 , g167 ); 
buf ( n169 , g168 ); 
buf ( n170 , g169 ); 
buf ( n171 , g170 ); 
buf ( n172 , g171 ); 
buf ( n173 , g172 ); 
buf ( n174 , g173 ); 
buf ( n175 , g174 ); 
buf ( n176 , g175 ); 
buf ( n177 , g176 ); 
buf ( n178 , g177 ); 
buf ( n179 , g178 ); 
buf ( n180 , g179 ); 
buf ( n181 , g180 ); 
buf ( n182 , g181 ); 
buf ( n183 , g182 ); 
buf ( n184 , g183 ); 
buf ( n185 , g184 ); 
buf ( n186 , g185 ); 
buf ( n187 , g186 ); 
buf ( n188 , g187 ); 
buf ( n189 , g188 ); 
buf ( n190 , g189 ); 
buf ( n191 , g190 ); 
buf ( n192 , g191 ); 
buf ( n193 , g192 ); 
buf ( n194 , g193 ); 
buf ( n195 , g194 ); 
buf ( n196 , g195 ); 
buf ( n197 , g196 ); 
buf ( n198 , g197 ); 
buf ( n199 , g198 ); 
buf ( n200 , g199 ); 
buf ( n201 , g200 ); 
buf ( n202 , g201 ); 
buf ( n203 , g202 ); 
buf ( n204 , g203 ); 
buf ( n205 , g204 ); 
buf ( n206 , g205 ); 
buf ( n207 , g206 ); 
buf ( g207 , n208 ); 
buf ( g208 , n209 ); 
buf ( g209 , n210 ); 
buf ( g210 , n211 ); 
buf ( g211 , n212 ); 
buf ( g212 , n213 ); 
buf ( g213 , n214 ); 
buf ( g214 , n215 ); 
buf ( g215 , n216 ); 
buf ( g216 , n217 ); 
buf ( g217 , n218 ); 
buf ( g218 , n219 ); 
buf ( g219 , n220 ); 
buf ( g220 , n221 ); 
buf ( g221 , n222 ); 
buf ( g222 , n223 ); 
buf ( g223 , n224 ); 
buf ( g224 , n225 ); 
buf ( g225 , n226 ); 
buf ( g226 , n227 ); 
buf ( g227 , n228 ); 
buf ( g228 , n229 ); 
buf ( g229 , n230 ); 
buf ( g230 , n231 ); 
buf ( n208 , n1747 ); 
buf ( n209 , n1338 ); 
buf ( n210 , n2162 ); 
buf ( n211 , n1460 ); 
buf ( n212 , n2207 ); 
buf ( n213 , n1595 ); 
buf ( n214 , n2252 ); 
buf ( n215 , n1651 ); 
buf ( n216 , n1699 ); 
buf ( n217 , n2300 ); 
buf ( n218 , n1200 ); 
buf ( n219 , n2118 ); 
buf ( n220 , n2344 ); 
buf ( n221 , n1853 ); 
buf ( n222 , n1898 ); 
buf ( n223 , n1952 ); 
buf ( n224 , n2002 ); 
buf ( n225 , n2050 ); 
buf ( n226 , n1805 ); 
buf ( n227 , n2419 ); 
buf ( n228 , n2826 ); 
buf ( n229 , n2922 ); 
buf ( n230 , n2873 ); 
buf ( n231 , n2723 ); 
not ( n237 , n96 ); 
or ( n238 , n237 , n2 , n67 ); 
not ( n239 , n3 ); 
nor ( n240 , n239 , n2 ); 
buf ( n241 , n240 ); 
not ( n242 , n241 ); 
not ( n243 , n242 ); 
not ( n244 , n243 ); 
not ( n245 , n244 ); 
not ( n246 , n245 ); 
not ( n247 , n246 ); 
not ( n248 , n247 ); 
not ( n249 , n248 ); 
not ( n250 , n7 ); 
nor ( n251 , n250 , n2 ); 
not ( n252 , n251 ); 
or ( n253 , n249 , n252 ); 
not ( n254 , n12 ); 
nor ( n255 , n254 , n2 ); 
not ( n256 , n255 ); 
not ( n257 , n2 ); 
nand ( n258 , n257 , n13 ); 
nand ( n259 , n256 , n258 ); 
not ( n260 , n14 ); 
nor ( n261 , n260 , n2 ); 
not ( n262 , n261 ); 
not ( n263 , n15 ); 
nor ( n264 , n263 , n2 ); 
not ( n265 , n264 ); 
nand ( n266 , n262 , n265 ); 
nor ( n267 , n259 , n266 ); 
not ( n268 , n267 ); 
not ( n269 , n2 ); 
nand ( n270 , n269 , n9 ); 
not ( n271 , n270 ); 
not ( n272 , n2 ); 
nand ( n273 , n272 , n8 ); 
not ( n274 , n2 ); 
nand ( n275 , n274 , n10 ); 
nand ( n276 , n273 , n275 ); 
not ( n277 , n2 ); 
nand ( n278 , n277 , n11 ); 
not ( n279 , n278 ); 
nor ( n280 , n268 , n271 , n276 , n279 ); 
not ( n281 , n2 ); 
nand ( n282 , n281 , n24 ); 
not ( n283 , n2 ); 
nand ( n284 , n283 , n25 ); 
nand ( n285 , n282 , n284 ); 
not ( n286 , n285 ); 
not ( n287 , n26 ); 
nor ( n288 , n287 , n2 ); 
not ( n289 , n27 ); 
nor ( n290 , n289 , n2 ); 
nor ( n291 , n288 , n290 ); 
nor ( n292 , n20 , n21 ); 
nor ( n293 , n292 , n2 ); 
not ( n294 , n293 ); 
not ( n295 , n2 ); 
nand ( n296 , n295 , n22 ); 
not ( n297 , n2 ); 
nand ( n298 , n297 , n23 ); 
and ( n299 , n296 , n298 ); 
nand ( n300 , n286 , n291 , n294 , n299 ); 
not ( n301 , n2 ); 
nand ( n302 , n301 , n16 ); 
not ( n303 , n2 ); 
nand ( n304 , n303 , n17 ); 
and ( n305 , n302 , n304 ); 
not ( n306 , n2 ); 
nand ( n307 , n306 , n18 ); 
not ( n308 , n2 ); 
nand ( n309 , n308 , n19 ); 
nand ( n310 , n307 , n309 ); 
not ( n311 , n310 ); 
nand ( n312 , n305 , n311 ); 
nor ( n313 , n300 , n312 ); 
not ( n314 , n28 ); 
nor ( n315 , n314 , n2 ); 
not ( n316 , n315 ); 
not ( n317 , n2 ); 
nand ( n318 , n317 , n29 ); 
nand ( n319 , n316 , n318 ); 
not ( n320 , n30 ); 
nor ( n321 , n320 , n2 ); 
not ( n322 , n321 ); 
not ( n323 , n2 ); 
nand ( n324 , n323 , n31 ); 
nand ( n325 , n322 , n324 ); 
nor ( n326 , n319 , n325 ); 
nand ( n327 , n313 , n326 ); 
not ( n328 , n327 ); 
and ( n329 , n280 , n328 ); 
not ( n330 , n329 ); 
or ( n331 , n251 , n330 ); 
and ( n332 , n251 , n330 ); 
not ( n333 , n242 ); 
buf ( n334 , n333 ); 
not ( n335 , n334 ); 
buf ( n336 , n335 ); 
nor ( n337 , n332 , n336 ); 
nand ( n338 , n331 , n337 ); 
nand ( n339 , n253 , n338 ); 
not ( n340 , n339 ); 
not ( n341 , n324 ); 
not ( n342 , n341 ); 
not ( n343 , n293 ); 
not ( n344 , n2 ); 
nand ( n345 , n344 , n22 ); 
buf ( n346 , n298 ); 
nand ( n347 , n343 , n345 , n346 ); 
not ( n348 , n347 ); 
not ( n349 , n291 ); 
not ( n350 , n349 ); 
nand ( n351 , n348 , n350 , n286 , n311 ); 
not ( n352 , n319 ); 
nand ( n353 , n352 , n305 ); 
nor ( n354 , n351 , n353 ); 
not ( n355 , n354 ); 
not ( n356 , n355 ); 
and ( n357 , n342 , n356 ); 
not ( n358 , n341 ); 
not ( n359 , n355 ); 
or ( n360 , n358 , n359 ); 
buf ( n361 , n243 ); 
nand ( n362 , n360 , n361 ); 
nor ( n363 , n357 , n362 ); 
buf ( n364 , n241 ); 
buf ( n365 , n364 ); 
not ( n366 , n341 ); 
nor ( n367 , n365 , n366 ); 
nor ( n368 , n363 , n367 ); 
not ( n369 , n304 ); 
not ( n370 , n369 ); 
nand ( n371 , n370 , n324 ); 
nor ( n372 , n371 , n319 ); 
not ( n373 , n290 ); 
and ( n374 , n373 , n296 ); 
not ( n375 , n23 ); 
nor ( n376 , n375 , n2 ); 
nor ( n377 , n293 , n376 ); 
nand ( n378 , n374 , n286 , n377 ); 
not ( n379 , n302 ); 
not ( n380 , n26 ); 
nor ( n381 , n380 , n2 ); 
nor ( n382 , n379 , n381 ); 
nand ( n383 , n382 , n311 ); 
nor ( n384 , n378 , n383 ); 
nand ( n385 , n372 , n384 ); 
not ( n386 , n321 ); 
not ( n387 , n386 ); 
nor ( n388 , n385 , n387 ); 
not ( n389 , n388 ); 
not ( n390 , n387 ); 
not ( n391 , n385 ); 
or ( n392 , n390 , n391 ); 
nand ( n393 , n392 , n365 ); 
not ( n394 , n393 ); 
and ( n395 , n389 , n394 ); 
not ( n396 , n364 ); 
and ( n397 , n396 , n387 ); 
nor ( n398 , n395 , n397 ); 
nand ( n399 , n368 , n398 ); 
not ( n400 , n244 ); 
not ( n401 , n307 ); 
not ( n402 , n401 ); 
not ( n403 , n402 ); 
not ( n404 , n403 ); 
or ( n405 , n400 , n404 ); 
not ( n406 , n402 ); 
not ( n407 , n300 ); 
not ( n408 , n407 ); 
or ( n409 , n406 , n408 ); 
not ( n410 , n401 ); 
not ( n411 , n300 ); 
or ( n412 , n410 , n411 ); 
nand ( n413 , n412 , n333 ); 
not ( n414 , n413 ); 
nand ( n415 , n409 , n414 ); 
nand ( n416 , n405 , n415 ); 
not ( n417 , n416 ); 
not ( n418 , n309 ); 
not ( n419 , n376 ); 
not ( n420 , n345 ); 
not ( n421 , n420 ); 
not ( n422 , n284 ); 
not ( n423 , n422 ); 
not ( n424 , n20 ); 
nor ( n425 , n424 , n2 ); 
not ( n426 , n21 ); 
nor ( n427 , n426 , n2 ); 
nor ( n428 , n425 , n427 ); 
nand ( n429 , n419 , n421 , n423 , n428 ); 
not ( n430 , n429 ); 
not ( n431 , n2 ); 
nand ( n432 , n431 , n24 ); 
and ( n433 , n307 , n432 ); 
not ( n434 , n433 ); 
nor ( n435 , n349 , n434 ); 
nand ( n436 , n430 , n435 ); 
not ( n437 , n436 ); 
not ( n438 , n437 ); 
or ( n439 , n418 , n438 ); 
not ( n440 , n19 ); 
nor ( n441 , n440 , n2 ); 
not ( n442 , n441 ); 
not ( n443 , n436 ); 
or ( n444 , n442 , n443 ); 
not ( n445 , n242 ); 
nand ( n446 , n444 , n445 ); 
not ( n447 , n446 ); 
nand ( n448 , n439 , n447 ); 
nand ( n449 , n242 , n441 ); 
nand ( n450 , n448 , n449 ); 
buf ( n451 , n379 ); 
not ( n452 , n451 ); 
not ( n453 , n351 ); 
or ( n454 , n452 , n453 ); 
nand ( n455 , n454 , n333 ); 
nor ( n456 , n451 , n351 ); 
or ( n457 , n455 , n456 ); 
not ( n458 , n451 ); 
or ( n459 , n365 , n458 ); 
nand ( n460 , n457 , n459 ); 
nor ( n461 , n450 , n460 ); 
nand ( n462 , n417 , n461 ); 
not ( n463 , n462 ); 
not ( n464 , n244 ); 
not ( n465 , n370 ); 
not ( n466 , n465 ); 
or ( n467 , n464 , n466 ); 
nor ( n468 , n370 , n384 ); 
not ( n469 , n468 ); 
nand ( n470 , n370 , n384 ); 
nand ( n471 , n469 , n470 , n361 ); 
nand ( n472 , n467 , n471 ); 
not ( n473 , n472 ); 
not ( n474 , n396 ); 
not ( n475 , n315 ); 
or ( n476 , n474 , n475 ); 
nor ( n477 , n316 , n313 ); 
not ( n478 , n477 ); 
nand ( n479 , n316 , n313 ); 
nand ( n480 , n478 , n479 , n365 ); 
nand ( n481 , n476 , n480 ); 
not ( n482 , n481 ); 
not ( n483 , n318 ); 
not ( n484 , n483 ); 
not ( n485 , n484 ); 
not ( n486 , n302 ); 
nor ( n487 , n486 , n369 ); 
nor ( n488 , n441 , n315 ); 
and ( n489 , n433 , n291 , n487 , n488 ); 
not ( n490 , n422 ); 
not ( n491 , n420 ); 
and ( n492 , n490 , n491 , n428 , n346 ); 
nand ( n493 , n489 , n492 ); 
not ( n494 , n493 ); 
not ( n495 , n494 ); 
or ( n496 , n485 , n495 ); 
nand ( n497 , n496 , n365 ); 
not ( n498 , n493 ); 
not ( n499 , n483 ); 
nor ( n500 , n498 , n499 ); 
or ( n501 , n497 , n500 ); 
or ( n502 , n361 , n499 ); 
nand ( n503 , n501 , n502 ); 
not ( n504 , n503 ); 
nand ( n505 , n473 , n482 , n504 ); 
not ( n506 , n505 ); 
nand ( n507 , n463 , n506 ); 
nor ( n508 , n399 , n507 ); 
not ( n509 , n265 ); 
not ( n510 , n509 ); 
nor ( n511 , n259 , n325 ); 
nand ( n512 , n354 , n511 ); 
not ( n513 , n512 ); 
or ( n514 , n510 , n513 ); 
nand ( n515 , n514 , n334 ); 
not ( n516 , n265 ); 
nor ( n517 , n516 , n512 ); 
or ( n518 , n515 , n517 ); 
not ( n519 , n516 ); 
or ( n520 , n245 , n519 ); 
nand ( n521 , n518 , n520 ); 
not ( n522 , n521 ); 
not ( n523 , n334 ); 
and ( n524 , n374 , n286 , n377 ); 
not ( n525 , n383 ); 
not ( n526 , n264 ); 
nand ( n527 , n526 , n386 ); 
nor ( n528 , n259 , n527 ); 
buf ( n529 , n528 ); 
and ( n530 , n524 , n372 , n525 , n529 ); 
not ( n531 , n530 ); 
not ( n532 , n262 ); 
and ( n533 , n531 , n532 ); 
not ( n534 , n524 ); 
not ( n535 , n372 ); 
nand ( n536 , n528 , n311 , n382 ); 
nor ( n537 , n534 , n535 , n536 ); 
and ( n538 , n537 , n262 ); 
nor ( n539 , n533 , n538 ); 
not ( n540 , n539 ); 
or ( n541 , n523 , n540 ); 
nand ( n542 , n396 , n261 ); 
nand ( n543 , n541 , n542 ); 
not ( n544 , n543 ); 
not ( n545 , n244 ); 
not ( n546 , n255 ); 
not ( n547 , n546 ); 
not ( n548 , n547 ); 
or ( n549 , n545 , n548 ); 
nor ( n550 , n547 , n327 ); 
not ( n551 , n550 ); 
nand ( n552 , n547 , n327 ); 
nand ( n553 , n551 , n552 , n365 ); 
nand ( n554 , n549 , n553 ); 
not ( n555 , n258 ); 
not ( n556 , n555 ); 
nand ( n557 , n546 , n318 ); 
nor ( n558 , n557 , n325 ); 
not ( n559 , n429 ); 
nand ( n560 , n559 , n489 , n558 ); 
nor ( n561 , n554 , t_0 ); 
nand ( n562 , n522 , n544 , n561 ); 
not ( n563 , n562 ); 
not ( n564 , n336 ); 
not ( n565 , n564 ); 
nand ( n566 , n267 , n328 ); 
and ( n567 , n566 , n270 ); 
not ( n568 , n566 ); 
and ( n569 , n568 , n271 ); 
nor ( n570 , n567 , n569 ); 
not ( n571 , n570 ); 
not ( n572 , n571 ); 
or ( n573 , n565 , n572 ); 
nand ( n574 , n335 , n271 ); 
nand ( n575 , n573 , n574 ); 
not ( n576 , n575 ); 
not ( n577 , n275 ); 
nand ( n578 , n336 , n577 ); 
not ( n579 , n275 ); 
and ( n580 , n273 , n270 , n278 , n262 ); 
nand ( n581 , n580 , n537 ); 
not ( n582 , n581 ); 
not ( n583 , n582 ); 
or ( n584 , n579 , n583 ); 
not ( n585 , n577 ); 
not ( n586 , n581 ); 
or ( n587 , n585 , n586 ); 
not ( n588 , n335 ); 
nand ( n589 , n587 , n588 ); 
not ( n590 , n589 ); 
nand ( n591 , n584 , n590 ); 
and ( n592 , n578 , n591 ); 
nand ( n593 , n576 , n592 ); 
not ( n594 , n377 ); 
nand ( n595 , n241 , n594 ); 
not ( n596 , n491 ); 
xor ( n597 , n595 , n596 ); 
not ( n598 , n425 ); 
not ( n599 , n598 ); 
not ( n600 , n599 ); 
nor ( n601 , n239 , n2 ); 
not ( n602 , n598 ); 
nand ( n603 , n601 , n602 ); 
not ( n604 , n21 ); 
nor ( n605 , n604 , n2 ); 
not ( n606 , n605 ); 
and ( n607 , n603 , n606 ); 
not ( n608 , n603 ); 
and ( n609 , n608 , n605 ); 
nor ( n610 , n607 , n609 ); 
not ( n611 , n610 ); 
not ( n612 , n294 ); 
nand ( n613 , n612 , n601 ); 
and ( n614 , n613 , n346 ); 
not ( n615 , n613 ); 
and ( n616 , n615 , n376 ); 
nor ( n617 , n614 , n616 ); 
not ( n618 , n617 ); 
and ( n619 , n597 , n600 , n611 , n618 ); 
not ( n620 , n619 ); 
not ( n621 , n620 ); 
not ( n622 , n286 ); 
not ( n623 , n348 ); 
or ( n624 , n622 , n623 ); 
nand ( n625 , n624 , n364 ); 
not ( n626 , n373 ); 
and ( n627 , n625 , n626 ); 
not ( n628 , n625 ); 
and ( n629 , n628 , n373 ); 
nor ( n630 , n627 , n629 ); 
not ( n631 , n396 ); 
not ( n632 , n381 ); 
or ( n633 , n631 , n632 ); 
not ( n634 , n381 ); 
not ( n635 , n634 ); 
not ( n636 , n524 ); 
or ( n637 , n635 , n636 ); 
not ( n638 , n381 ); 
not ( n639 , n378 ); 
or ( n640 , n638 , n639 ); 
nand ( n641 , n640 , n445 ); 
not ( n642 , n641 ); 
nand ( n643 , n637 , n642 ); 
nand ( n644 , n633 , n643 ); 
not ( n645 , n644 ); 
not ( n646 , n294 ); 
not ( n647 , n299 ); 
or ( n648 , n646 , n647 ); 
nand ( n649 , n648 , n241 ); 
not ( n650 , n490 ); 
and ( n651 , n649 , n650 ); 
not ( n652 , n649 ); 
and ( n653 , n652 , n490 ); 
nor ( n654 , n651 , n653 ); 
not ( n655 , n654 ); 
not ( n656 , n492 ); 
nand ( n657 , n656 , n364 ); 
buf ( n658 , n432 ); 
and ( n659 , n657 , n658 ); 
not ( n660 , n657 ); 
not ( n661 , n658 ); 
and ( n662 , n660 , n661 ); 
nor ( n663 , n659 , n662 ); 
nor ( n664 , n655 , n663 ); 
and ( n665 , n630 , n645 , n664 ); 
not ( n666 , n665 ); 
not ( n667 , n246 ); 
not ( n668 , n279 ); 
or ( n669 , n667 , n668 ); 
nor ( n670 , n271 , n266 ); 
nand ( n671 , n670 , n556 ); 
nor ( n672 , n560 , n671 ); 
nor ( n673 , n278 , n672 ); 
not ( n674 , n673 ); 
not ( n675 , n671 ); 
not ( n676 , n560 ); 
nand ( n677 , n278 , n675 , n676 ); 
nand ( n678 , n674 , n677 , n588 ); 
nand ( n679 , n669 , n678 ); 
nor ( n680 , n666 , n679 ); 
not ( n681 , n273 ); 
not ( n682 , n355 ); 
not ( n683 , n682 ); 
nand ( n684 , n670 , n278 , n511 ); 
nor ( n685 , n683 , n684 ); 
not ( n686 , n685 ); 
or ( n687 , n681 , n686 ); 
not ( n688 , n273 ); 
not ( n689 , n688 ); 
not ( n690 , n685 ); 
not ( n691 , n690 ); 
or ( n692 , n689 , n691 ); 
not ( n693 , n246 ); 
nand ( n694 , n692 , n693 ); 
not ( n695 , n694 ); 
nand ( n696 , n687 , n695 ); 
not ( n697 , n696 ); 
nor ( n698 , n245 , n273 ); 
nor ( n699 , n697 , n698 ); 
nand ( n700 , n621 , n680 , n699 ); 
nor ( n701 , n593 , n700 ); 
nand ( n702 , n508 , n563 , n701 ); 
not ( n703 , n2 ); 
nand ( n704 , n703 , n1 ); 
not ( n705 , n704 ); 
not ( n706 , n2 ); 
nand ( n707 , n706 , n32 ); 
not ( n708 , n707 ); 
nor ( n709 , n705 , n708 ); 
not ( n710 , n2 ); 
nand ( n711 , n710 , n33 ); 
not ( n712 , n2 ); 
nand ( n713 , n712 , n4 ); 
and ( n714 , n580 , n529 ); 
nor ( n715 , n251 , n577 ); 
not ( n716 , n2 ); 
nand ( n717 , n716 , n5 ); 
not ( n718 , n2 ); 
nand ( n719 , n718 , n6 ); 
nand ( n720 , n717 , n719 ); 
nor ( n721 , n720 , n385 ); 
and ( n722 , n713 , n714 , n715 , n721 ); 
and ( n723 , n709 , n711 , n588 , n722 ); 
buf ( n724 , n723 ); 
nand ( n725 , n702 , n724 ); 
and ( n726 , n340 , n725 ); 
and ( n727 , n336 , n719 ); 
not ( n728 , n336 ); 
not ( n729 , n276 ); 
not ( n730 , n251 ); 
nand ( n731 , n729 , n730 , n278 ); 
not ( n732 , n731 ); 
and ( n733 , n305 , n488 ); 
and ( n734 , n733 , n558 , n675 ); 
buf ( n735 , n437 ); 
nand ( n736 , n732 , n734 , n735 ); 
nand ( n737 , n719 , n736 ); 
and ( n738 , n728 , n737 ); 
nor ( n739 , n727 , n738 ); 
nor ( n740 , n736 , n335 , n719 ); 
nor ( n741 , n739 , n740 ); 
not ( n742 , n741 ); 
nor ( n743 , n340 , n725 ); 
not ( n744 , n743 ); 
not ( n745 , n744 ); 
or ( n746 , n742 , n745 ); 
not ( n747 , n741 ); 
nand ( n748 , n747 , n743 ); 
nand ( n749 , n746 , n748 ); 
nor ( n750 , n726 , n749 ); 
nor ( n751 , n246 , n717 ); 
not ( n752 , n751 ); 
not ( n753 , n276 ); 
and ( n754 , n719 , n730 ); 
nand ( n755 , n753 , n685 , n754 ); 
not ( n756 , n755 ); 
not ( n757 , n756 ); 
or ( n758 , n752 , n757 ); 
not ( n759 , n717 ); 
nor ( n760 , n759 , n588 ); 
not ( n761 , n760 ); 
not ( n762 , n717 ); 
not ( n763 , n755 ); 
or ( n764 , n762 , n763 ); 
nand ( n765 , n764 , n247 ); 
nand ( n766 , n761 , n765 ); 
nand ( n767 , n758 , n766 ); 
not ( n768 , n767 ); 
buf ( n769 , n768 ); 
buf ( n770 , n769 ); 
not ( n771 , n770 ); 
not ( n772 , n748 ); 
and ( n773 , n771 , n772 ); 
and ( n774 , n770 , n748 ); 
nor ( n775 , n773 , n774 ); 
and ( n776 , n750 , n744 , n775 ); 
buf ( n777 , n776 ); 
not ( n778 , n777 ); 
not ( n779 , n778 ); 
not ( n780 , n460 ); 
not ( n781 , n780 ); 
not ( n782 , n542 ); 
nor ( n783 , n679 , n782 ); 
not ( n784 , n574 ); 
nor ( n785 , n698 , n784 ); 
not ( n786 , n539 ); 
not ( n787 , n786 ); 
not ( n788 , n570 ); 
or ( n789 , n787 , n788 ); 
nand ( n790 , n789 , n564 ); 
and ( n791 , n696 , n783 , n785 , n790 ); 
buf ( n792 , n521 ); 
not ( n793 , n792 ); 
not ( n794 , n398 ); 
not ( n795 , n794 ); 
nand ( n796 , n793 , n795 , n561 ); 
not ( n797 , n796 ); 
and ( n798 , n791 , n797 ); 
and ( n799 , n592 , n340 ); 
buf ( n800 , n482 ); 
not ( n801 , n800 ); 
not ( n802 , n504 ); 
nor ( n803 , n801 , n802 ); 
not ( n804 , n472 ); 
buf ( n805 , n804 ); 
not ( n806 , n368 ); 
not ( n807 , n806 ); 
nand ( n808 , n803 , n805 , n807 ); 
not ( n809 , n808 ); 
and ( n810 , n630 , n619 , n664 ); 
not ( n811 , n810 ); 
not ( n812 , n644 ); 
not ( n813 , n812 ); 
not ( n814 , n416 ); 
not ( n815 , n814 ); 
nor ( n816 , n813 , n815 ); 
buf ( n817 , n461 ); 
nand ( n818 , n816 , n817 ); 
nor ( n819 , n811 , n818 ); 
nand ( n820 , n809 , n768 , n741 , n819 ); 
not ( n821 , n820 ); 
nand ( n822 , n798 , n799 , n821 ); 
and ( n823 , n724 , n822 ); 
not ( n824 , n713 ); 
nand ( n825 , n824 , n248 ); 
not ( n826 , n714 ); 
nand ( n827 , n715 , n721 ); 
nor ( n828 , n826 , n827 ); 
or ( n829 , n713 , n828 ); 
not ( n830 , n722 ); 
nand ( n831 , n829 , n830 , n564 ); 
and ( n832 , n825 , n831 ); 
not ( n833 , n832 ); 
nor ( n834 , n823 , n833 ); 
not ( n835 , n834 ); 
nand ( n836 , n835 , 1'b1 ); 
not ( n837 , n836 ); 
and ( n838 , n713 , n717 ); 
nand ( n839 , n754 , n838 , n329 ); 
nor ( n840 , n705 , n839 ); 
not ( n841 , n705 ); 
not ( n842 , n839 ); 
or ( n843 , n841 , n842 ); 
nand ( n844 , n843 , n564 ); 
or ( n845 , n840 , n844 ); 
not ( n846 , n248 ); 
or ( n847 , n846 , n704 ); 
nand ( n848 , n845 , n847 ); 
not ( n849 , n848 ); 
and ( n850 , 1'b1 , n849 ); 
nor ( n851 , n850 , 1'b0 ); 
not ( n852 , n851 ); 
nand ( n853 , n837 , n852 ); 
not ( n854 , n853 ); 
not ( n855 , n854 ); 
not ( n856 , n855 ); 
nand ( n857 , n781 , n856 ); 
not ( n858 , n836 ); 
nand ( n859 , n858 , n851 ); 
buf ( n860 , n859 ); 
not ( n861 , n860 ); 
not ( n862 , n2 ); 
nand ( n863 , n43 , n862 ); 
nor ( n864 , n863 , n780 ); 
not ( n865 , n864 ); 
nand ( n866 , n863 , n780 ); 
nand ( n867 , n865 , n866 ); 
not ( n868 , n417 ); 
or ( n869 , n46 , n868 ); 
not ( n870 , n44 ); 
nor ( n871 , n870 , n2 ); 
or ( n872 , n871 , n450 ); 
and ( n873 , n869 , n872 ); 
not ( n874 , n873 ); 
not ( n875 , n2 ); 
nand ( n876 , n875 , n45 ); 
nand ( n877 , n876 , n812 ); 
not ( n878 , n877 ); 
not ( n879 , n630 ); 
nor ( n880 , n879 , n40 ); 
nor ( n881 , n878 , n880 ); 
not ( n882 , n881 ); 
not ( n883 , n2 ); 
nand ( n884 , n883 , n42 ); 
nand ( n885 , n884 , n654 ); 
not ( n886 , n885 ); 
not ( n887 , n39 ); 
not ( n888 , n663 ); 
nand ( n889 , n887 , n888 ); 
not ( n890 , n889 ); 
nor ( n891 , n886 , n890 ); 
not ( n892 , n891 ); 
not ( n893 , n2 ); 
nand ( n894 , n893 , n36 ); 
not ( n895 , n894 ); 
and ( n896 , n895 , n610 ); 
not ( n897 , n896 ); 
not ( n898 , n2 ); 
nand ( n899 , n898 , n38 ); 
not ( n900 , n899 ); 
and ( n901 , n599 , n900 ); 
nand ( n902 , n894 , n611 ); 
nand ( n903 , n901 , n902 ); 
nand ( n904 , n897 , n903 ); 
not ( n905 , n904 ); 
not ( n906 , n2 ); 
nand ( n907 , n906 , n37 ); 
not ( n908 , n617 ); 
nand ( n909 , n907 , n908 ); 
not ( n910 , n2 ); 
nand ( n911 , n910 , n41 ); 
nand ( n912 , n911 , n597 ); 
and ( n913 , n909 , n912 ); 
not ( n914 , n913 ); 
or ( n915 , n905 , n914 ); 
nor ( n916 , n911 , n597 ); 
not ( n917 , n916 ); 
nor ( n918 , n907 , n908 ); 
nand ( n919 , n918 , n912 ); 
nand ( n920 , n917 , n919 ); 
not ( n921 , n920 ); 
nand ( n922 , n915 , n921 ); 
not ( n923 , n922 ); 
or ( n924 , n892 , n923 ); 
nand ( n925 , n39 , n663 ); 
nor ( n926 , n884 , n654 ); 
nand ( n927 , n926 , n889 ); 
nand ( n928 , n925 , n927 ); 
not ( n929 , n928 ); 
nand ( n930 , n924 , n929 ); 
not ( n931 , n930 ); 
or ( n932 , n882 , n931 ); 
nand ( n933 , n40 , n879 ); 
not ( n934 , n933 ); 
and ( n935 , n934 , n877 ); 
nor ( n936 , n876 , n645 ); 
nor ( n937 , n935 , n936 ); 
nand ( n938 , n932 , n937 ); 
not ( n939 , n938 ); 
or ( n940 , n874 , n939 ); 
not ( n941 , n417 ); 
buf ( n942 , n941 ); 
and ( n943 , n46 , n942 ); 
and ( n944 , n943 , n872 ); 
and ( n945 , n871 , n450 ); 
nor ( n946 , n944 , n945 ); 
nand ( n947 , n940 , n946 ); 
not ( n948 , n947 ); 
xor ( n949 , n867 , n948 ); 
nand ( n950 , n861 , n949 ); 
not ( n951 , n95 ); 
nor ( n952 , n951 , n2 ); 
nand ( n953 , n852 , n836 ); 
not ( n954 , n953 ); 
not ( n955 , n954 ); 
not ( n956 , n955 ); 
nand ( n957 , n952 , n956 ); 
nand ( n958 , n836 , n851 ); 
buf ( n959 , n958 ); 
not ( n960 , n959 ); 
nand ( n961 , n59 , n862 ); 
nor ( n962 , n961 , n780 ); 
not ( n963 , n962 ); 
nand ( n964 , n780 , n961 ); 
nand ( n965 , n963 , n964 ); 
not ( n966 , n965 ); 
nand ( n967 , n62 , n862 ); 
nand ( n968 , n967 , n814 ); 
not ( n969 , n2 ); 
nand ( n970 , n969 , n60 ); 
not ( n971 , n450 ); 
nand ( n972 , n970 , n971 ); 
buf ( n973 , n972 ); 
and ( n974 , n968 , n973 ); 
not ( n975 , n974 ); 
not ( n976 , n2 ); 
nand ( n977 , n976 , n56 ); 
nand ( n978 , n977 , n630 ); 
not ( n979 , n2 ); 
nand ( n980 , n979 , n61 ); 
nand ( n981 , n980 , n645 ); 
and ( n982 , n978 , n981 ); 
not ( n983 , n982 ); 
not ( n984 , n2 ); 
nand ( n985 , n984 , n58 ); 
nand ( n986 , n985 , n654 ); 
not ( n987 , n986 ); 
not ( n988 , n663 ); 
not ( n989 , n2 ); 
nand ( n990 , n989 , n55 ); 
nand ( n991 , n988 , n990 ); 
not ( n992 , n991 ); 
nor ( n993 , n987 , n992 ); 
not ( n994 , n993 ); 
not ( n995 , n2 ); 
nand ( n996 , n995 , n52 ); 
not ( n997 , n996 ); 
and ( n998 , n997 , n610 ); 
not ( n999 , n998 ); 
not ( n1000 , n2 ); 
nand ( n1001 , n1000 , n54 ); 
not ( n1002 , n1001 ); 
and ( n1003 , n599 , n1002 ); 
nand ( n1004 , n996 , n611 ); 
nand ( n1005 , n1003 , n1004 ); 
nand ( n1006 , n999 , n1005 ); 
not ( n1007 , n1006 ); 
not ( n1008 , n617 ); 
not ( n1009 , n2 ); 
nand ( n1010 , n1009 , n53 ); 
nand ( n1011 , n1008 , n1010 ); 
not ( n1012 , n2 ); 
nand ( n1013 , n1012 , n57 ); 
nand ( n1014 , n1013 , n597 ); 
and ( n1015 , n1011 , n1014 ); 
not ( n1016 , n1015 ); 
or ( n1017 , n1007 , n1016 ); 
nor ( n1018 , n1013 , n597 ); 
not ( n1019 , n1018 ); 
not ( n1020 , n617 ); 
nor ( n1021 , n1010 , n1020 ); 
nand ( n1022 , n1021 , n1014 ); 
nand ( n1023 , n1019 , n1022 ); 
not ( n1024 , n1023 ); 
nand ( n1025 , n1017 , n1024 ); 
not ( n1026 , n1025 ); 
or ( n1027 , n994 , n1026 ); 
not ( n1028 , n663 ); 
nor ( n1029 , n990 , n1028 ); 
not ( n1030 , n1029 ); 
nor ( n1031 , n985 , n654 ); 
nand ( n1032 , n1031 , n991 ); 
nand ( n1033 , n1030 , n1032 ); 
not ( n1034 , n1033 ); 
nand ( n1035 , n1027 , n1034 ); 
not ( n1036 , n1035 ); 
or ( n1037 , n983 , n1036 ); 
nor ( n1038 , n977 , n630 ); 
buf ( n1039 , n1038 ); 
and ( n1040 , n1039 , n981 ); 
not ( n1041 , n980 ); 
and ( n1042 , n1041 , n813 ); 
nor ( n1043 , n1040 , n1042 ); 
nand ( n1044 , n1037 , n1043 ); 
not ( n1045 , n1044 ); 
or ( n1046 , n975 , n1045 ); 
not ( n1047 , n967 ); 
and ( n1048 , n1047 , n941 ); 
and ( n1049 , n1048 , n973 ); 
nor ( n1050 , n971 , n970 ); 
buf ( n1051 , n1050 ); 
nor ( n1052 , n1049 , n1051 ); 
nand ( n1053 , n1046 , n1052 ); 
nand ( n1054 , n966 , n1053 ); 
not ( n1055 , n1053 ); 
nand ( n1056 , n965 , n1055 ); 
nand ( n1057 , n960 , n1054 , n1056 ); 
nand ( n1058 , n857 , n950 , n957 , n1057 ); 
not ( n1059 , n1058 ); 
not ( n1060 , n723 ); 
not ( n1061 , n562 ); 
nor ( n1062 , n399 , n462 , n505 ); 
nand ( n1063 , n1061 , n1062 , n665 ); 
not ( n1064 , n1063 ); 
or ( n1065 , n1060 , n1064 ); 
nand ( n1066 , n620 , n723 ); 
nand ( n1067 , n1065 , n1066 ); 
buf ( n1068 , n1067 ); 
and ( n1069 , n1068 , n575 ); 
not ( n1070 , n1068 ); 
and ( n1071 , n1070 , n576 ); 
nor ( n1072 , n1069 , n1071 ); 
buf ( n1073 , n1072 ); 
nand ( n1074 , n1067 , n575 ); 
not ( n1075 , n1074 ); 
not ( n1076 , n679 ); 
not ( n1077 , n1076 ); 
nand ( n1078 , n1075 , n1077 ); 
buf ( n1079 , n699 ); 
nor ( n1080 , n1078 , n1079 ); 
not ( n1081 , n592 ); 
and ( n1082 , n1080 , n1081 ); 
not ( n1083 , n1080 ); 
and ( n1084 , n1083 , n592 ); 
nor ( n1085 , n1082 , n1084 ); 
nor ( n1086 , n1073 , n1085 ); 
not ( n1087 , n1086 ); 
not ( n1088 , n1087 ); 
not ( n1089 , n1076 ); 
not ( n1090 , n1089 ); 
not ( n1091 , n1075 ); 
not ( n1092 , n1091 ); 
or ( n1093 , n1090 , n1092 ); 
or ( n1094 , n1089 , n1091 ); 
nand ( n1095 , n1093 , n1094 ); 
buf ( n1096 , n1095 ); 
not ( n1097 , n1078 ); 
not ( n1098 , n1079 ); 
and ( n1099 , n1097 , n1098 ); 
not ( n1100 , n1097 ); 
and ( n1101 , n1100 , n1079 ); 
nor ( n1102 , n1099 , n1101 ); 
not ( n1103 , n1102 ); 
nor ( n1104 , n1096 , n1103 ); 
nand ( n1105 , n1088 , n1104 ); 
not ( n1106 , n1087 ); 
nor ( n1107 , n1096 , n1102 ); 
nand ( n1108 , n1106 , n1107 ); 
nand ( n1109 , n1105 , n1108 ); 
not ( n1110 , n1085 ); 
nand ( n1111 , n1110 , n1073 ); 
not ( n1112 , n1111 ); 
nand ( n1113 , n1112 , n1107 ); 
not ( n1114 , n1111 ); 
nand ( n1115 , n1114 , n1104 ); 
nand ( n1116 , n1113 , n1115 ); 
nor ( n1117 , n1109 , n1116 ); 
not ( n1118 , n1102 ); 
nand ( n1119 , n1118 , n1096 ); 
not ( n1120 , n1119 ); 
nand ( n1121 , n1096 , n1102 , n1086 ); 
not ( n1122 , n1121 ); 
or ( n1123 , n1120 , n1122 ); 
nand ( n1124 , n1111 , n1087 ); 
nand ( n1125 , n1123 , n1124 ); 
not ( n1126 , n1107 ); 
nand ( n1127 , n1073 , n1085 ); 
not ( n1128 , n1127 ); 
not ( n1129 , n1128 ); 
or ( n1130 , n1126 , n1129 ); 
not ( n1131 , n1119 ); 
not ( n1132 , n1073 ); 
nand ( n1133 , n1132 , n1085 ); 
nand ( n1134 , n1127 , n1133 ); 
nand ( n1135 , n1131 , n1134 ); 
nand ( n1136 , n1130 , n1135 ); 
not ( n1137 , n1136 ); 
and ( n1138 , n1117 , n1125 , n1137 ); 
not ( n1139 , n1107 ); 
not ( n1140 , n1133 ); 
not ( n1141 , n1140 ); 
or ( n1142 , n1139 , n1141 ); 
not ( n1143 , n1111 ); 
nand ( n1144 , n1143 , n1102 , n1096 ); 
nand ( n1145 , n1142 , n1144 ); 
not ( n1146 , n1145 ); 
nand ( n1147 , n1138 , n1146 ); 
not ( n1148 , n1147 ); 
or ( n1149 , n1059 , n1148 ); 
not ( n1150 , n1104 ); 
not ( n1151 , n1140 ); 
or ( n1152 , n1150 , n1151 ); 
not ( n1153 , n1073 ); 
not ( n1154 , n1096 ); 
nand ( n1155 , n1153 , n1154 ); 
not ( n1156 , n1110 ); 
nand ( n1157 , n1155 , n1102 , n1156 ); 
nand ( n1158 , n1152 , n1157 ); 
buf ( n1159 , n1158 ); 
nand ( n1160 , n952 , n1159 ); 
nand ( n1161 , n1149 , n1160 ); 
not ( n1162 , n1161 ); 
or ( n1163 , n779 , n1162 ); 
nor ( n1164 , n808 , n818 ); 
and ( n1165 , n797 , n1164 ); 
buf ( n1166 , n810 ); 
buf ( n1167 , n791 ); 
nand ( n1168 , n1165 , n1166 , n1167 ); 
nand ( n1169 , n724 , n1168 ); 
and ( n1170 , n1169 , n592 ); 
not ( n1171 , n1169 ); 
and ( n1172 , n1171 , n1081 ); 
or ( n1173 , n1170 , n1172 ); 
not ( n1174 , n1173 ); 
not ( n1175 , n1174 ); 
nand ( n1176 , n1163 , n1175 ); 
not ( n1177 , n781 ); 
not ( n1178 , n1177 ); 
not ( n1179 , n955 ); 
not ( n1180 , n1179 ); 
not ( n1181 , n1180 ); 
and ( n1182 , n1178 , n1181 ); 
not ( n1183 , n950 ); 
nor ( n1184 , n1182 , n1183 ); 
not ( n1185 , n1057 ); 
not ( n1186 , n857 ); 
nor ( n1187 , n1185 , n1186 ); 
and ( n1188 , n1184 , n1187 ); 
not ( n1189 , n777 ); 
nor ( n1190 , n1188 , n1189 ); 
nor ( n1191 , n1176 , n1190 ); 
buf ( n1192 , n1173 ); 
not ( n1193 , n1192 ); 
not ( n1194 , n1193 ); 
not ( n1195 , n1058 ); 
not ( n1196 , n1195 ); 
or ( n1197 , n1194 , n1196 ); 
nand ( n1198 , n1197 , n67 ); 
or ( n1199 , n1191 , n1198 ); 
nand ( n1200 , n238 , n1199 ); 
not ( n1201 , n72 ); 
or ( n1202 , n1201 , n2 , n67 ); 
not ( n1203 , n778 ); 
not ( n1204 , n71 ); 
nor ( n1205 , n1204 , n2 ); 
buf ( n1206 , n954 ); 
nand ( n1207 , n1205 , n1206 ); 
not ( n1208 , n860 ); 
nand ( n1209 , n69 , n862 ); 
buf ( n1210 , n554 ); 
not ( n1211 , n1210 ); 
buf ( n1212 , n1211 ); 
buf ( n1213 , n1212 ); 
nor ( n1214 , n1209 , n1213 ); 
not ( n1215 , n1214 ); 
nand ( n1216 , n1209 , n1211 ); 
nand ( n1217 , n1215 , n1216 ); 
nand ( n1218 , n47 , n862 ); 
nand ( n1219 , n1218 , n805 ); 
and ( n1220 , n864 , n1219 ); 
nor ( n1221 , n1218 , n804 ); 
nor ( n1222 , n1220 , n1221 ); 
and ( n1223 , n866 , n1219 ); 
nand ( n1224 , n1223 , n947 ); 
nand ( n1225 , n1222 , n1224 ); 
nand ( n1226 , n48 , n862 ); 
nand ( n1227 , n1226 , n800 ); 
nand ( n1228 , n49 , n862 ); 
not ( n1229 , n802 ); 
nand ( n1230 , n1228 , n1229 ); 
nand ( n1231 , n1225 , n1227 , n1230 ); 
nand ( n1232 , n50 , n862 ); 
not ( n1233 , n806 ); 
nand ( n1234 , n1232 , n1233 ); 
nand ( n1235 , n35 , n862 ); 
not ( n1236 , n794 ); 
nand ( n1237 , n1235 , n1236 ); 
nand ( n1238 , n1234 , n1237 ); 
or ( n1239 , n1231 , n1238 ); 
not ( n1240 , n1235 ); 
not ( n1241 , n795 ); 
nand ( n1242 , n1240 , n1241 ); 
nand ( n1243 , n1239 , n1242 ); 
nor ( n1244 , n1232 , n1233 ); 
not ( n1245 , n1244 ); 
not ( n1246 , n1237 ); 
or ( n1247 , n1245 , n1246 ); 
nor ( n1248 , n1226 , n800 ); 
and ( n1249 , n1248 , n1230 ); 
not ( n1250 , n802 ); 
nor ( n1251 , n1250 , n1228 ); 
nor ( n1252 , n1249 , n1251 ); 
or ( n1253 , n1238 , n1252 ); 
nand ( n1254 , n1247 , n1253 ); 
nor ( n1255 , n1243 , n1254 ); 
nand ( n1256 , n1217 , n1255 ); 
not ( n1257 , n1217 ); 
not ( n1258 , n1255 ); 
nand ( n1259 , n1257 , n1258 ); 
nand ( n1260 , n1208 , n1256 , n1259 ); 
not ( n1261 , n1213 ); 
not ( n1262 , n855 ); 
nand ( n1263 , n1261 , n1262 ); 
not ( n1264 , n959 ); 
nand ( n1265 , n70 , n862 ); 
not ( n1266 , n1210 ); 
nand ( n1267 , n1265 , n1266 ); 
not ( n1268 , n1267 ); 
nor ( n1269 , n1265 , n1212 ); 
nor ( n1270 , n1268 , n1269 ); 
nand ( n1271 , n63 , n862 ); 
nand ( n1272 , n1271 , n805 ); 
and ( n1273 , n962 , n1272 ); 
nor ( n1274 , n1271 , n804 ); 
nor ( n1275 , n1273 , n1274 ); 
and ( n1276 , n964 , n1272 ); 
nand ( n1277 , n1276 , n1053 ); 
nand ( n1278 , n1275 , n1277 ); 
nand ( n1279 , n64 , n862 ); 
nand ( n1280 , n1279 , n800 ); 
nand ( n1281 , n65 , n862 ); 
nand ( n1282 , n1281 , n1250 ); 
nand ( n1283 , n1278 , n1280 , n1282 ); 
nand ( n1284 , n66 , n862 ); 
not ( n1285 , n806 ); 
nand ( n1286 , n1284 , n1285 ); 
nand ( n1287 , n51 , n862 ); 
nand ( n1288 , n1287 , n398 ); 
nand ( n1289 , n1286 , n1288 ); 
or ( n1290 , n1283 , n1289 ); 
not ( n1291 , n1287 ); 
nand ( n1292 , n1291 , n1241 ); 
not ( n1293 , n1292 ); 
not ( n1294 , n1293 ); 
nand ( n1295 , n1290 , n1294 ); 
nor ( n1296 , n1284 , n1233 ); 
not ( n1297 , n1296 ); 
not ( n1298 , n1288 ); 
or ( n1299 , n1297 , n1298 ); 
nor ( n1300 , n1279 , n800 ); 
and ( n1301 , n1300 , n1282 ); 
nor ( n1302 , n1281 , n1250 ); 
nor ( n1303 , n1301 , n1302 ); 
or ( n1304 , n1289 , n1303 ); 
nand ( n1305 , n1299 , n1304 ); 
nor ( n1306 , n1295 , n1305 ); 
not ( n1307 , n1306 ); 
nand ( n1308 , n1270 , n1307 ); 
not ( n1309 , n1270 ); 
nand ( n1310 , n1309 , n1306 ); 
nand ( n1311 , n1264 , n1308 , n1310 ); 
nand ( n1312 , n1207 , n1260 , n1263 , n1311 ); 
not ( n1313 , n1312 ); 
nand ( n1314 , n1138 , n1146 ); 
not ( n1315 , n1314 ); 
or ( n1316 , n1313 , n1315 ); 
nand ( n1317 , n1205 , n1159 ); 
nand ( n1318 , n1316 , n1317 ); 
not ( n1319 , n1318 ); 
or ( n1320 , n1203 , n1319 ); 
not ( n1321 , n1192 ); 
not ( n1322 , n1321 ); 
nand ( n1323 , n1320 , n1322 ); 
nand ( n1324 , n1261 , n1179 ); 
and ( n1325 , n1324 , n1260 ); 
not ( n1326 , n1311 ); 
not ( n1327 , n1263 ); 
nor ( n1328 , n1326 , n1327 ); 
and ( n1329 , n1325 , n1328 ); 
nor ( n1330 , n1329 , n1189 ); 
nor ( n1331 , n1323 , n1330 ); 
not ( n1332 , n1193 ); 
not ( n1333 , n1312 ); 
not ( n1334 , n1333 ); 
or ( n1335 , n1332 , n1334 ); 
nand ( n1336 , n1335 , n67 ); 
or ( n1337 , n1331 , n1336 ); 
nand ( n1338 , n1202 , n1337 ); 
not ( n1339 , n67 ); 
nand ( n1340 , n76 , n862 , n1339 ); 
not ( n1341 , n1250 ); 
buf ( n1342 , n1206 ); 
and ( n1343 , n1341 , n1342 ); 
not ( n1344 , n860 ); 
not ( n1345 , n1251 ); 
nand ( n1346 , n1345 , n1230 ); 
nand ( n1347 , n1219 , n1227 ); 
and ( n1348 , n945 , n866 ); 
nor ( n1349 , n1348 , n864 ); 
or ( n1350 , n1347 , n1349 ); 
and ( n1351 , n1221 , n1227 ); 
nor ( n1352 , n1351 , n1248 ); 
nand ( n1353 , n1350 , n1352 ); 
and ( n1354 , n936 , n869 ); 
nor ( n1355 , n1354 , n943 ); 
and ( n1356 , n877 , n869 ); 
or ( n1357 , n925 , n880 ); 
nand ( n1358 , n1357 , n933 ); 
not ( n1359 , n1358 ); 
nor ( n1360 , n890 , n880 ); 
not ( n1361 , n918 ); 
nand ( n1362 , n896 , n909 ); 
nand ( n1363 , n1361 , n1362 ); 
not ( n1364 , n909 ); 
nor ( n1365 , n1364 , n903 ); 
or ( n1366 , n1363 , n1365 ); 
and ( n1367 , n912 , n885 ); 
nand ( n1368 , n1366 , n1367 ); 
and ( n1369 , n916 , n885 ); 
nor ( n1370 , n1369 , n926 ); 
nand ( n1371 , n1368 , n1370 ); 
nand ( n1372 , n1360 , n1371 ); 
nand ( n1373 , n1359 , n1372 ); 
nand ( n1374 , n1356 , n1373 ); 
nand ( n1375 , n1355 , n1374 ); 
not ( n1376 , n1375 ); 
nand ( n1377 , n872 , n866 ); 
buf ( n1378 , n1377 ); 
buf ( n1379 , n1378 ); 
nor ( n1380 , n1376 , n1379 , n1347 ); 
nor ( n1381 , n1353 , n1380 ); 
nand ( n1382 , n1346 , n1381 ); 
or ( n1383 , n1346 , n1381 ); 
nand ( n1384 , n1344 , n1382 , n1383 ); 
not ( n1385 , n1384 ); 
nor ( n1386 , n1343 , n1385 ); 
not ( n1387 , n959 ); 
not ( n1388 , n1302 ); 
nand ( n1389 , n1388 , n1282 ); 
nand ( n1390 , n1272 , n1280 ); 
and ( n1391 , n1051 , n964 ); 
nor ( n1392 , n1391 , n962 ); 
or ( n1393 , n1390 , n1392 ); 
and ( n1394 , n1274 , n1280 ); 
nor ( n1395 , n1394 , n1300 ); 
nand ( n1396 , n1393 , n1395 ); 
and ( n1397 , n981 , n968 ); 
not ( n1398 , n1397 ); 
and ( n1399 , n1014 , n986 ); 
not ( n1400 , n1399 ); 
and ( n1401 , n998 , n1011 ); 
nor ( n1402 , n1401 , n1021 ); 
nor ( n1403 , n1400 , n1402 ); 
not ( n1404 , n1011 ); 
nor ( n1405 , n1404 , n1005 ); 
not ( n1406 , n1405 ); 
not ( n1407 , n1399 ); 
or ( n1408 , n1406 , n1407 ); 
and ( n1409 , n1018 , n986 ); 
nor ( n1410 , n1409 , n1031 ); 
nand ( n1411 , n1408 , n1410 ); 
nor ( n1412 , n1403 , n1411 ); 
nand ( n1413 , n991 , n978 ); 
or ( n1414 , n1412 , n1413 ); 
and ( n1415 , n1029 , n978 ); 
nor ( n1416 , n1415 , n1038 ); 
nand ( n1417 , n1414 , n1416 ); 
not ( n1418 , n1417 ); 
or ( n1419 , n1398 , n1418 ); 
and ( n1420 , n1042 , n968 ); 
nor ( n1421 , n1420 , n1048 ); 
nand ( n1422 , n1419 , n1421 ); 
not ( n1423 , n1422 ); 
nand ( n1424 , n964 , n972 ); 
nor ( n1425 , n1423 , n1424 , n1390 ); 
nor ( n1426 , n1396 , n1425 ); 
nand ( n1427 , n1389 , n1426 ); 
not ( n1428 , n1389 ); 
not ( n1429 , n1426 ); 
nand ( n1430 , n1428 , n1429 ); 
nand ( n1431 , n1387 , n1427 , n1430 ); 
not ( n1432 , n1431 ); 
nand ( n1433 , n1341 , n1262 ); 
not ( n1434 , n1433 ); 
nor ( n1435 , n1432 , n1434 ); 
and ( n1436 , n1386 , n1435 ); 
not ( n1437 , n777 ); 
nor ( n1438 , n1436 , n1437 ); 
not ( n1439 , n1438 ); 
not ( n1440 , n777 ); 
not ( n1441 , n75 ); 
nor ( n1442 , n1441 , n2 ); 
nand ( n1443 , n1442 , n1206 ); 
nand ( n1444 , n1443 , n1384 , n1433 , n1431 ); 
not ( n1445 , n1444 ); 
and ( n1446 , n1108 , n1113 , n1105 , n1115 ); 
nand ( n1447 , n1446 , n1146 , n1125 , n1137 ); 
not ( n1448 , n1447 ); 
or ( n1449 , n1445 , n1448 ); 
nand ( n1450 , n1442 , n1159 ); 
nand ( n1451 , n1449 , n1450 ); 
nand ( n1452 , n1440 , n1451 ); 
not ( n1453 , n1192 ); 
not ( n1454 , n1453 ); 
nand ( n1455 , n1439 , n1452 , n1454 ); 
not ( n1456 , n1444 ); 
and ( n1457 , n1321 , n1456 ); 
nor ( n1458 , n1457 , n1339 ); 
nand ( n1459 , n1455 , n1458 ); 
nand ( n1460 , n1340 , n1459 ); 
not ( n1461 , n86 ); 
or ( n1462 , n1461 , n2 , n67 ); 
not ( n1463 , n860 ); 
nand ( n1464 , n79 , n862 ); 
not ( n1465 , n543 ); 
not ( n1466 , n1465 ); 
and ( n1467 , n1464 , n1466 ); 
not ( n1468 , n1464 ); 
and ( n1469 , n1468 , n1465 ); 
nor ( n1470 , n1467 , n1469 ); 
nand ( n1471 , n1237 , n1216 ); 
nand ( n1472 , n80 , n862 ); 
buf ( n1473 , t_0 ); 
not ( n1474 , n1473 ); 
nand ( n1475 , n1472 , n1474 ); 
nand ( n1476 , n81 , n862 ); 
not ( n1477 , n792 ); 
nand ( n1478 , n1476 , n1477 ); 
nand ( n1479 , n1475 , n1478 ); 
nor ( n1480 , n1471 , n1479 ); 
or ( n1481 , n1355 , n1378 ); 
nand ( n1482 , n1481 , n1349 ); 
not ( n1483 , n1377 ); 
nand ( n1484 , n1483 , n1356 ); 
not ( n1485 , n1365 ); 
not ( n1486 , n1363 ); 
nand ( n1487 , n1485 , n1486 ); 
nand ( n1488 , n1487 , n1367 , n1360 ); 
not ( n1489 , n1358 ); 
not ( n1490 , n1370 ); 
nand ( n1491 , n1490 , n1360 ); 
and ( n1492 , n1488 , n1489 , n1491 ); 
nor ( n1493 , n1484 , n1492 ); 
nor ( n1494 , n1482 , n1493 ); 
nand ( n1495 , n1230 , n1234 ); 
nor ( n1496 , n1494 , n1347 , n1495 ); 
and ( n1497 , n1480 , n1496 ); 
not ( n1498 , n1242 ); 
and ( n1499 , n1498 , n1216 ); 
nor ( n1500 , n1499 , n1214 ); 
or ( n1501 , n1500 , n1479 ); 
or ( n1502 , n1495 , n1352 ); 
and ( n1503 , n1234 , n1251 ); 
nor ( n1504 , n1503 , n1244 ); 
nand ( n1505 , n1502 , n1504 ); 
nand ( n1506 , n1480 , n1505 ); 
nand ( n1507 , n1501 , n1506 ); 
buf ( n1508 , n1477 ); 
or ( n1509 , n1476 , n1508 ); 
buf ( n1510 , n1474 ); 
nor ( n1511 , n1472 , n1510 ); 
nand ( n1512 , n1511 , n1478 ); 
nand ( n1513 , n1509 , n1512 ); 
nor ( n1514 , n1497 , n1507 , n1513 ); 
nand ( n1515 , n1470 , n1514 ); 
or ( n1516 , n1470 , n1514 ); 
nand ( n1517 , n1463 , n1515 , n1516 ); 
not ( n1518 , n82 ); 
nor ( n1519 , n1518 , n2 ); 
not ( n1520 , n955 ); 
nand ( n1521 , n1519 , n1520 ); 
not ( n1522 , n855 ); 
nand ( n1523 , n1522 , n1466 ); 
not ( n1524 , n959 ); 
nand ( n1525 , n83 , n862 ); 
xor ( n1526 , n1525 , n1465 ); 
not ( n1527 , n1526 ); 
nand ( n1528 , n84 , n862 ); 
buf ( n1529 , n1510 ); 
nor ( n1530 , n1528 , n1529 ); 
not ( n1531 , n85 ); 
nor ( n1532 , n1531 , n2 ); 
or ( n1533 , n1532 , n792 ); 
and ( n1534 , n1530 , n1533 ); 
not ( n1535 , n1508 ); 
and ( n1536 , n1532 , n1535 ); 
nor ( n1537 , n1534 , n1536 ); 
nand ( n1538 , n1288 , n1267 ); 
not ( n1539 , n1473 ); 
nand ( n1540 , n1528 , n1539 ); 
nand ( n1541 , n1540 , n1533 ); 
nor ( n1542 , n1538 , n1541 ); 
or ( n1543 , n1421 , n1424 ); 
nand ( n1544 , n1543 , n1392 ); 
or ( n1545 , n1413 , n1410 ); 
not ( n1546 , n1413 ); 
not ( n1547 , n1405 ); 
nand ( n1548 , n1547 , n1402 ); 
nand ( n1549 , n1546 , n1399 , n1548 ); 
nand ( n1550 , n1545 , n1549 , n1416 ); 
not ( n1551 , n1424 ); 
and ( n1552 , n1550 , n1397 , n1551 ); 
nor ( n1553 , n1544 , n1552 ); 
nand ( n1554 , n1282 , n1286 ); 
nor ( n1555 , n1553 , n1390 , n1554 ); 
and ( n1556 , n1542 , n1555 ); 
and ( n1557 , n1293 , n1267 ); 
nor ( n1558 , n1557 , n1269 ); 
or ( n1559 , n1541 , n1558 ); 
or ( n1560 , n1554 , n1395 ); 
and ( n1561 , n1286 , n1302 ); 
nor ( n1562 , n1561 , n1296 ); 
nand ( n1563 , n1560 , n1562 ); 
nand ( n1564 , n1542 , n1563 ); 
nand ( n1565 , n1559 , n1564 ); 
nor ( n1566 , n1556 , n1565 ); 
nand ( n1567 , n1537 , n1566 ); 
not ( n1568 , n1567 ); 
nand ( n1569 , n1527 , n1568 ); 
nand ( n1570 , n1526 , n1567 ); 
nand ( n1571 , n1524 , n1569 , n1570 ); 
nand ( n1572 , n1517 , n1521 , n1523 , n1571 ); 
and ( n1573 , n1321 , n1572 ); 
not ( n1574 , n1321 ); 
not ( n1575 , n777 ); 
not ( n1576 , n1575 ); 
not ( n1577 , n1447 ); 
not ( n1578 , n1572 ); 
or ( n1579 , n1577 , n1578 ); 
nand ( n1580 , n1159 , n1519 ); 
nand ( n1581 , n1579 , n1580 ); 
not ( n1582 , n1581 ); 
or ( n1583 , n1576 , n1582 ); 
not ( n1584 , n1466 ); 
not ( n1585 , n1342 ); 
or ( n1586 , n1584 , n1585 ); 
nand ( n1587 , n1586 , n1523 ); 
nand ( n1588 , n1517 , n1571 ); 
or ( n1589 , n1587 , n1588 ); 
nand ( n1590 , n1589 , n777 ); 
nand ( n1591 , n1583 , n1590 ); 
and ( n1592 , n1574 , n1591 ); 
nor ( n1593 , n1573 , n1592 ); 
or ( n1594 , n1593 , n1339 ); 
nand ( n1595 , n1462 , n1594 ); 
not ( n1596 , n90 ); 
or ( n1597 , n1596 , n2 , n67 ); 
not ( n1598 , n777 ); 
not ( n1599 , n1598 ); 
not ( n1600 , n1285 ); 
not ( n1601 , n855 ); 
nand ( n1602 , n1600 , n1601 ); 
not ( n1603 , n860 ); 
not ( n1604 , n1244 ); 
nand ( n1605 , n1604 , n1234 ); 
nand ( n1606 , n1252 , n1231 ); 
not ( n1607 , n1606 ); 
nand ( n1608 , n1605 , n1607 ); 
not ( n1609 , n1605 ); 
nand ( n1610 , n1609 , n1606 ); 
nand ( n1611 , n1603 , n1608 , n1610 ); 
not ( n1612 , n89 ); 
nor ( n1613 , n1612 , n2 ); 
nand ( n1614 , n1613 , n1206 ); 
not ( n1615 , n959 ); 
not ( n1616 , n1296 ); 
nand ( n1617 , n1616 , n1286 ); 
nand ( n1618 , n1303 , n1283 ); 
not ( n1619 , n1618 ); 
nand ( n1620 , n1617 , n1619 ); 
not ( n1621 , n1617 ); 
nand ( n1622 , n1621 , n1618 ); 
nand ( n1623 , n1615 , n1620 , n1622 ); 
nand ( n1624 , n1602 , n1611 , n1614 , n1623 ); 
not ( n1625 , n1624 ); 
nand ( n1626 , n1138 , n1146 ); 
not ( n1627 , n1626 ); 
or ( n1628 , n1625 , n1627 ); 
nand ( n1629 , n1613 , n1159 ); 
nand ( n1630 , n1628 , n1629 ); 
not ( n1631 , n1630 ); 
or ( n1632 , n1599 , n1631 ); 
not ( n1633 , n1321 ); 
nand ( n1634 , n1632 , n1633 ); 
not ( n1635 , n955 ); 
buf ( n1636 , n1635 ); 
nand ( n1637 , n1600 , n1636 ); 
and ( n1638 , n1637 , n1611 ); 
not ( n1639 , n1623 ); 
not ( n1640 , n1602 ); 
nor ( n1641 , n1639 , n1640 ); 
and ( n1642 , n1638 , n1641 ); 
nor ( n1643 , n1642 , n1189 ); 
nor ( n1644 , n1634 , n1643 ); 
not ( n1645 , n1193 ); 
not ( n1646 , n1624 ); 
not ( n1647 , n1646 ); 
or ( n1648 , n1645 , n1647 ); 
nand ( n1649 , n1648 , n67 ); 
or ( n1650 , n1644 , n1649 ); 
nand ( n1651 , n1597 , n1650 ); 
not ( n1652 , n92 ); 
or ( n1653 , n1652 , n2 , n67 ); 
not ( n1654 , n778 ); 
not ( n1655 , n959 ); 
not ( n1656 , n1274 ); 
nand ( n1657 , n1656 , n1272 ); 
not ( n1658 , n1657 ); 
not ( n1659 , n1553 ); 
nand ( n1660 , n1658 , n1659 ); 
nand ( n1661 , n1657 , n1553 ); 
nand ( n1662 , n1655 , n1660 , n1661 ); 
not ( n1663 , n860 ); 
not ( n1664 , n1221 ); 
nand ( n1665 , n1664 , n1219 ); 
nand ( n1666 , n1665 , n1494 ); 
not ( n1667 , n1665 ); 
not ( n1668 , n1494 ); 
nand ( n1669 , n1667 , n1668 ); 
nand ( n1670 , n1663 , n1666 , n1669 ); 
not ( n1671 , n805 ); 
nand ( n1672 , n1671 , n1262 ); 
not ( n1673 , n91 ); 
nor ( n1674 , n1673 , n2 ); 
nand ( n1675 , n1674 , n1635 ); 
nand ( n1676 , n1662 , n1670 , n1672 , n1675 ); 
not ( n1677 , n1676 ); 
not ( n1678 , n1314 ); 
or ( n1679 , n1677 , n1678 ); 
nand ( n1680 , n1674 , n1159 ); 
nand ( n1681 , n1679 , n1680 ); 
not ( n1682 , n1681 ); 
or ( n1683 , n1654 , n1682 ); 
nand ( n1684 , n1683 , n1322 ); 
nand ( n1685 , n1671 , n1179 ); 
and ( n1686 , n1685 , n1670 ); 
not ( n1687 , n1662 ); 
not ( n1688 , n1672 ); 
nor ( n1689 , n1687 , n1688 ); 
and ( n1690 , n1686 , n1689 ); 
nor ( n1691 , n1690 , n1189 ); 
nor ( n1692 , n1684 , n1691 ); 
not ( n1693 , n1193 ); 
not ( n1694 , n1676 ); 
not ( n1695 , n1694 ); 
or ( n1696 , n1693 , n1695 ); 
nand ( n1697 , n1696 , n67 ); 
or ( n1698 , n1692 , n1697 ); 
nand ( n1699 , n1653 , n1698 ); 
not ( n1700 , n68 ); 
or ( n1701 , n1700 , n2 , n67 ); 
not ( n1702 , n777 ); 
not ( n1703 , n1702 ); 
nand ( n1704 , n1241 , n1601 ); 
not ( n1705 , n860 ); 
nand ( n1706 , n1242 , n1237 ); 
nor ( n1707 , n1505 , n1496 ); 
nand ( n1708 , n1706 , n1707 ); 
not ( n1709 , n1706 ); 
not ( n1710 , n1707 ); 
nand ( n1711 , n1709 , n1710 ); 
nand ( n1712 , n1705 , n1708 , n1711 ); 
not ( n1713 , n959 ); 
nand ( n1714 , n1294 , n1288 ); 
not ( n1715 , n1714 ); 
nor ( n1716 , n1563 , n1555 ); 
not ( n1717 , n1716 ); 
nand ( n1718 , n1715 , n1717 ); 
nand ( n1719 , n1714 , n1716 ); 
nand ( n1720 , n1713 , n1718 , n1719 ); 
not ( n1721 , n34 ); 
nor ( n1722 , n1721 , n2 ); 
nand ( n1723 , n1722 , n1206 ); 
nand ( n1724 , n1704 , n1712 , n1720 , n1723 ); 
not ( n1725 , n1724 ); 
not ( n1726 , n1626 ); 
or ( n1727 , n1725 , n1726 ); 
nand ( n1728 , n1722 , n1159 ); 
nand ( n1729 , n1727 , n1728 ); 
not ( n1730 , n1729 ); 
or ( n1731 , n1703 , n1730 ); 
nand ( n1732 , n1731 , n1633 ); 
nand ( n1733 , n1241 , n1636 ); 
and ( n1734 , n1733 , n1712 ); 
not ( n1735 , n1720 ); 
not ( n1736 , n1704 ); 
nor ( n1737 , n1735 , n1736 ); 
and ( n1738 , n1734 , n1737 ); 
nor ( n1739 , n1738 , n1189 ); 
nor ( n1740 , n1732 , n1739 ); 
not ( n1741 , n1321 ); 
not ( n1742 , n1724 ); 
not ( n1743 , n1742 ); 
or ( n1744 , n1741 , n1743 ); 
nand ( n1745 , n1744 , n67 ); 
or ( n1746 , n1740 , n1745 ); 
nand ( n1747 , n1701 , n1746 ); 
nand ( n1748 , n112 , n862 , n1339 ); 
not ( n1749 , n777 ); 
not ( n1750 , n853 ); 
nand ( n1751 , n1750 , n610 ); 
not ( n1752 , n958 ); 
not ( n1753 , n1003 ); 
not ( n1754 , n1004 ); 
nor ( n1755 , n1754 , n998 ); 
xnor ( n1756 , n1753 , n1755 ); 
nand ( n1757 , n1752 , n1756 ); 
nand ( n1758 , n1751 , n1757 ); 
not ( n1759 , n610 ); 
not ( n1760 , n1179 ); 
or ( n1761 , n1759 , n1760 ); 
not ( n1762 , n859 ); 
not ( n1763 , n901 ); 
not ( n1764 , n902 ); 
nor ( n1765 , n1764 , n896 ); 
not ( n1766 , n1765 ); 
nand ( n1767 , n1763 , n1766 ); 
not ( n1768 , n1763 ); 
nand ( n1769 , n1768 , n1765 ); 
nand ( n1770 , n1762 , n1767 , n1769 ); 
nand ( n1771 , n1761 , n1770 ); 
nor ( n1772 , n1758 , n1771 ); 
nor ( n1773 , n1749 , n1772 ); 
not ( n1774 , n1773 ); 
nand ( n1775 , n1113 , n1105 ); 
not ( n1776 , n1775 ); 
nand ( n1777 , n111 , n954 ); 
nand ( n1778 , n1757 , n1770 , n1751 , n1777 ); 
not ( n1779 , n1778 ); 
or ( n1780 , n1776 , n1779 ); 
nand ( n1781 , n111 , n1158 ); 
nand ( n1782 , n1780 , n1781 ); 
buf ( n1783 , n1108 ); 
not ( n1784 , n1778 ); 
nor ( n1785 , n1783 , n1784 ); 
nor ( n1786 , n1782 , n1785 ); 
not ( n1787 , n1786 ); 
not ( n1788 , n1115 ); 
nor ( n1789 , n1788 , n1145 ); 
nand ( n1790 , n1789 , n1125 , n1137 ); 
nand ( n1791 , n1790 , n1778 ); 
not ( n1792 , n1791 ); 
or ( n1793 , n1787 , n1792 ); 
not ( n1794 , n777 ); 
nand ( n1795 , n1793 , n1794 ); 
not ( n1796 , n1192 ); 
not ( n1797 , n1796 ); 
nand ( n1798 , n1774 , n1795 , n1797 ); 
not ( n1799 , n1784 ); 
not ( n1800 , n1174 ); 
or ( n1801 , n1799 , n1800 ); 
nand ( n1802 , n1801 , n67 ); 
not ( n1803 , n1802 ); 
nand ( n1804 , n1798 , n1803 ); 
nand ( n1805 , n1748 , n1804 ); 
nand ( n1806 , n102 , n862 , n1339 ); 
not ( n1807 , n800 ); 
nand ( n1808 , n1807 , n856 ); 
not ( n1809 , n1808 ); 
not ( n1810 , n959 ); 
not ( n1811 , n1300 ); 
nand ( n1812 , n1811 , n1280 ); 
not ( n1813 , n1812 ); 
nand ( n1814 , n1813 , n1278 ); 
not ( n1815 , n1278 ); 
nand ( n1816 , n1812 , n1815 ); 
nand ( n1817 , n1810 , n1814 , n1816 ); 
not ( n1818 , n1817 ); 
nor ( n1819 , n1809 , n1818 ); 
and ( n1820 , n1807 , n1179 ); 
not ( n1821 , n860 ); 
not ( n1822 , n1248 ); 
nand ( n1823 , n1822 , n1227 ); 
not ( n1824 , n1225 ); 
nand ( n1825 , n1823 , n1824 ); 
not ( n1826 , n1823 ); 
nand ( n1827 , n1826 , n1225 ); 
nand ( n1828 , n1821 , n1825 , n1827 ); 
not ( n1829 , n1828 ); 
nor ( n1830 , n1820 , n1829 ); 
and ( n1831 , n1819 , n1830 ); 
not ( n1832 , n777 ); 
nor ( n1833 , n1831 , n1832 ); 
not ( n1834 , n1833 ); 
not ( n1835 , n101 ); 
nor ( n1836 , n1835 , n2 ); 
nand ( n1837 , n1836 , n1206 ); 
nand ( n1838 , n1837 , n1828 , n1808 , n1817 ); 
not ( n1839 , n1838 ); 
nand ( n1840 , n1125 , n1137 ); 
not ( n1841 , n1840 ); 
nand ( n1842 , n1841 , n1146 , n1446 ); 
not ( n1843 , n1842 ); 
or ( n1844 , n1839 , n1843 ); 
nand ( n1845 , n1836 , n1159 ); 
nand ( n1846 , n1844 , n1845 ); 
nand ( n1847 , n1440 , n1846 ); 
nand ( n1848 , n1834 , n1847 , n1454 ); 
not ( n1849 , n1838 ); 
and ( n1850 , n1796 , n1849 ); 
nor ( n1851 , n1850 , n1339 ); 
nand ( n1852 , n1848 , n1851 ); 
nand ( n1853 , n1806 , n1852 ); 
nand ( n1854 , n104 , n862 , n1339 ); 
not ( n1855 , n600 ); 
not ( n1856 , n1855 ); 
not ( n1857 , n1856 ); 
nand ( n1858 , n1857 , n854 ); 
not ( n1859 , n958 ); 
nand ( n1860 , n1856 , n1001 ); 
nand ( n1861 , n1859 , n1860 , n1753 ); 
nand ( n1862 , n1858 , n1861 ); 
not ( n1863 , n1857 ); 
not ( n1864 , n1179 ); 
or ( n1865 , n1863 , n1864 ); 
not ( n1866 , n859 ); 
nand ( n1867 , n1856 , n899 ); 
nand ( n1868 , n1866 , n1867 , n1763 ); 
nand ( n1869 , n1865 , n1868 ); 
nor ( n1870 , n1862 , n1869 ); 
nor ( n1871 , n1575 , n1870 ); 
not ( n1872 , n1871 ); 
not ( n1873 , n1775 ); 
not ( n1874 , n103 ); 
nor ( n1875 , n1874 , n2 ); 
nand ( n1876 , n1875 , n954 ); 
nand ( n1877 , n1868 , n1861 , n1876 , n1858 ); 
not ( n1878 , n1877 ); 
or ( n1879 , n1873 , n1878 ); 
nand ( n1880 , n1875 , n1158 ); 
nand ( n1881 , n1879 , n1880 ); 
not ( n1882 , n1877 ); 
nor ( n1883 , n1783 , n1882 ); 
nor ( n1884 , n1881 , n1883 ); 
not ( n1885 , n1884 ); 
nand ( n1886 , n1790 , n1877 ); 
not ( n1887 , n1886 ); 
or ( n1888 , n1885 , n1887 ); 
nand ( n1889 , n1888 , n1794 ); 
buf ( n1890 , n1192 ); 
nand ( n1891 , n1872 , n1889 , n1890 ); 
not ( n1892 , n1882 ); 
not ( n1893 , n1174 ); 
or ( n1894 , n1892 , n1893 ); 
nand ( n1895 , n1894 , n67 ); 
not ( n1896 , n1895 ); 
nand ( n1897 , n1891 , n1896 ); 
nand ( n1898 , n1854 , n1897 ); 
not ( n1899 , n1339 ); 
not ( n1900 , n106 ); 
nor ( n1901 , n1900 , n2 ); 
not ( n1902 , n1901 ); 
or ( n1903 , n1899 , n1902 ); 
nand ( n1904 , n655 , n1750 ); 
not ( n1905 , n958 ); 
nor ( n1906 , n987 , n1031 ); 
not ( n1907 , n1906 ); 
not ( n1908 , n1025 ); 
nand ( n1909 , n1907 , n1908 ); 
nand ( n1910 , n1906 , n1025 ); 
nand ( n1911 , n1905 , n1909 , n1910 ); 
nand ( n1912 , n1904 , n1911 ); 
not ( n1913 , n655 ); 
not ( n1914 , n1342 ); 
or ( n1915 , n1913 , n1914 ); 
not ( n1916 , n859 ); 
nor ( n1917 , n886 , n926 ); 
not ( n1918 , n1917 ); 
not ( n1919 , n922 ); 
nand ( n1920 , n1918 , n1919 ); 
nand ( n1921 , n1917 , n922 ); 
nand ( n1922 , n1916 , n1920 , n1921 ); 
nand ( n1923 , n1915 , n1922 ); 
nor ( n1924 , n1912 , n1923 ); 
nor ( n1925 , n1749 , n1924 ); 
not ( n1926 , n1925 ); 
not ( n1927 , n1321 ); 
not ( n1928 , n1775 ); 
not ( n1929 , n105 ); 
nor ( n1930 , n1929 , n2 ); 
nand ( n1931 , n1930 , n954 ); 
nand ( n1932 , n1904 , n1922 , n1931 , n1911 ); 
not ( n1933 , n1932 ); 
or ( n1934 , n1928 , n1933 ); 
nand ( n1935 , n1930 , n1158 ); 
nand ( n1936 , n1934 , n1935 ); 
not ( n1937 , n1932 ); 
nor ( n1938 , n1783 , n1937 ); 
nor ( n1939 , n1936 , n1938 ); 
not ( n1940 , n1939 ); 
nand ( n1941 , n1790 , n1932 ); 
not ( n1942 , n1941 ); 
or ( n1943 , n1940 , n1942 ); 
nand ( n1944 , n1943 , n1794 ); 
nand ( n1945 , n1926 , n1927 , n1944 ); 
not ( n1946 , n1937 ); 
not ( n1947 , n1174 ); 
or ( n1948 , n1946 , n1947 ); 
nand ( n1949 , n1948 , n67 ); 
not ( n1950 , n1949 ); 
nand ( n1951 , n1945 , n1950 ); 
nand ( n1952 , n1903 , n1951 ); 
not ( n1953 , n1339 ); 
not ( n1954 , n108 ); 
nor ( n1955 , n1954 , n2 ); 
not ( n1956 , n1955 ); 
or ( n1957 , n1953 , n1956 ); 
not ( n1958 , n597 ); 
nand ( n1959 , n1958 , n1750 ); 
not ( n1960 , n958 ); 
not ( n1961 , n1014 ); 
nor ( n1962 , n1961 , n1018 ); 
xor ( n1963 , n1962 , n1548 ); 
nand ( n1964 , n1960 , n1963 ); 
nand ( n1965 , n1959 , n1964 ); 
not ( n1966 , n1958 ); 
not ( n1967 , n1635 ); 
or ( n1968 , n1966 , n1967 ); 
not ( n1969 , n859 ); 
not ( n1970 , n912 ); 
nor ( n1971 , n1970 , n916 ); 
xor ( n1972 , n1971 , n1487 ); 
nand ( n1973 , n1969 , n1972 ); 
nand ( n1974 , n1968 , n1973 ); 
nor ( n1975 , n1965 , n1974 ); 
nor ( n1976 , n1749 , n1975 ); 
not ( n1977 , n1976 ); 
not ( n1978 , n1775 ); 
nand ( n1979 , n107 , n954 ); 
nand ( n1980 , n1964 , n1979 , n1959 , n1973 ); 
not ( n1981 , n1980 ); 
or ( n1982 , n1978 , n1981 ); 
nand ( n1983 , n107 , n1158 ); 
nand ( n1984 , n1982 , n1983 ); 
not ( n1985 , n1980 ); 
nor ( n1986 , n1783 , n1985 ); 
nor ( n1987 , n1984 , n1986 ); 
not ( n1988 , n1987 ); 
nand ( n1989 , n1790 , n1980 ); 
not ( n1990 , n1989 ); 
or ( n1991 , n1988 , n1990 ); 
nand ( n1992 , n1991 , n1598 ); 
not ( n1993 , n1192 ); 
not ( n1994 , n1993 ); 
nand ( n1995 , n1977 , n1992 , n1994 ); 
not ( n1996 , n1985 ); 
not ( n1997 , n1174 ); 
or ( n1998 , n1996 , n1997 ); 
nand ( n1999 , n1998 , n67 ); 
not ( n2000 , n1999 ); 
nand ( n2001 , n1995 , n2000 ); 
nand ( n2002 , n1957 , n2001 ); 
not ( n2003 , n110 ); 
not ( n2004 , n1339 ); 
or ( n2005 , n2003 , n2004 ); 
not ( n2006 , n618 ); 
buf ( n2007 , n2006 ); 
not ( n2008 , n2007 ); 
not ( n2009 , n1342 ); 
or ( n2010 , n2008 , n2009 ); 
not ( n2011 , n859 ); 
not ( n2012 , n909 ); 
nor ( n2013 , n2012 , n918 ); 
or ( n2014 , n904 , n2013 ); 
nand ( n2015 , n904 , n2013 ); 
nand ( n2016 , n2011 , n2014 , n2015 ); 
nand ( n2017 , n2010 , n2016 ); 
nand ( n2018 , n1750 , n2007 ); 
not ( n2019 , n958 ); 
not ( n2020 , n1011 ); 
nor ( n2021 , n2020 , n1021 ); 
xor ( n2022 , n1006 , n2021 ); 
nand ( n2023 , n2019 , n2022 ); 
nand ( n2024 , n2018 , n2023 ); 
nor ( n2025 , n2017 , n2024 ); 
nor ( n2026 , n2025 , n1749 ); 
not ( n2027 , n2026 ); 
not ( n2028 , n1775 ); 
nand ( n2029 , n954 , n109 ); 
nand ( n2030 , n2023 , n2016 , n2018 , n2029 ); 
not ( n2031 , n2030 ); 
or ( n2032 , n2028 , n2031 ); 
nand ( n2033 , n109 , n1158 ); 
nand ( n2034 , n2032 , n2033 ); 
not ( n2035 , n2030 ); 
nor ( n2036 , n2035 , n1783 ); 
nor ( n2037 , n2034 , n2036 ); 
not ( n2038 , n2037 ); 
nand ( n2039 , n1790 , n2030 ); 
not ( n2040 , n2039 ); 
or ( n2041 , n2038 , n2040 ); 
nand ( n2042 , n2041 , n1598 ); 
nand ( n2043 , n2027 , n1797 , n2042 ); 
not ( n2044 , n2035 ); 
not ( n2045 , n1174 ); 
or ( n2046 , n2044 , n2045 ); 
nand ( n2047 , n2046 , n67 ); 
not ( n2048 , n2047 ); 
nand ( n2049 , n2043 , n2048 ); 
nand ( n2050 , n2005 , n2049 ); 
not ( n2051 , n98 ); 
or ( n2052 , n2051 , n2 , n67 ); 
not ( n2053 , n1702 ); 
not ( n2054 , n97 ); 
nor ( n2055 , n2054 , n2 ); 
nand ( n2056 , n2055 , n1206 ); 
not ( n2057 , n860 ); 
not ( n2058 , n1511 ); 
nand ( n2059 , n2058 , n1475 ); 
nor ( n2060 , n1495 , n1471 ); 
and ( n2061 , n2060 , n1353 ); 
not ( n2062 , n2060 ); 
not ( n2063 , n1380 ); 
or ( n2064 , n2062 , n2063 ); 
nand ( n2065 , n2064 , n1500 ); 
nor ( n2066 , n1471 , n1504 ); 
nor ( n2067 , n2061 , n2065 , n2066 ); 
nand ( n2068 , n2059 , n2067 ); 
not ( n2069 , n2059 ); 
not ( n2070 , n2067 ); 
nand ( n2071 , n2069 , n2070 ); 
nand ( n2072 , n2057 , n2068 , n2071 ); 
not ( n2073 , n1529 ); 
nand ( n2074 , n2073 , n1262 ); 
not ( n2075 , n959 ); 
not ( n2076 , n1530 ); 
nand ( n2077 , n2076 , n1540 ); 
not ( n2078 , n2077 ); 
nor ( n2079 , n1554 , n1538 ); 
and ( n2080 , n2079 , n1396 ); 
not ( n2081 , n2079 ); 
not ( n2082 , n1425 ); 
or ( n2083 , n2081 , n2082 ); 
nand ( n2084 , n2083 , n1558 ); 
nor ( n2085 , n1538 , n1562 ); 
nor ( n2086 , n2080 , n2084 , n2085 ); 
not ( n2087 , n2086 ); 
nand ( n2088 , n2078 , n2087 ); 
nand ( n2089 , n2077 , n2086 ); 
nand ( n2090 , n2075 , n2088 , n2089 ); 
nand ( n2091 , n2056 , n2072 , n2074 , n2090 ); 
not ( n2092 , n2091 ); 
not ( n2093 , n1147 ); 
or ( n2094 , n2092 , n2093 ); 
nand ( n2095 , n2055 , n1159 ); 
nand ( n2096 , n2094 , n2095 ); 
not ( n2097 , n2096 ); 
or ( n2098 , n2053 , n2097 ); 
nand ( n2099 , n2098 , n1927 ); 
not ( n2100 , n2073 ); 
not ( n2101 , n2100 ); 
not ( n2102 , n1180 ); 
and ( n2103 , n2101 , n2102 ); 
not ( n2104 , n2072 ); 
nor ( n2105 , n2103 , n2104 ); 
not ( n2106 , n2074 ); 
not ( n2107 , n2090 ); 
nor ( n2108 , n2106 , n2107 ); 
and ( n2109 , n2105 , n2108 ); 
nor ( n2110 , n2109 , n1189 ); 
nor ( n2111 , n2099 , n2110 ); 
not ( n2112 , n1453 ); 
not ( n2113 , n2091 ); 
not ( n2114 , n2113 ); 
or ( n2115 , n2112 , n2114 ); 
nand ( n2116 , n2115 , n67 ); 
or ( n2117 , n2111 , n2116 ); 
nand ( n2118 , n2052 , n2117 ); 
nand ( n2119 , n879 , n1636 ); 
not ( n2120 , n860 ); 
nor ( n2121 , n880 , n934 ); 
xor ( n2122 , n2121 , n930 ); 
nand ( n2123 , n2120 , n2122 ); 
and ( n2124 , n2119 , n2123 ); 
not ( n2125 , n959 ); 
not ( n2126 , n1039 ); 
nand ( n2127 , n2126 , n978 ); 
not ( n2128 , n2127 ); 
and ( n2129 , n1035 , n2128 ); 
not ( n2130 , n1035 ); 
and ( n2131 , n2130 , n2127 ); 
nor ( n2132 , n2129 , n2131 ); 
nand ( n2133 , n2125 , n2132 ); 
not ( n2134 , n2133 ); 
nand ( n2135 , n879 , n1601 ); 
not ( n2136 , n2135 ); 
nor ( n2137 , n2134 , n2136 ); 
and ( n2138 , n2124 , n2137 ); 
nor ( n2139 , n2138 , n1189 ); 
not ( n2140 , n1702 ); 
not ( n2141 , n73 ); 
nor ( n2142 , n2141 , n2 ); 
nand ( n2143 , n2142 , n956 ); 
nand ( n2144 , n2143 , n2123 , n2135 , n2133 ); 
not ( n2145 , n2144 ); 
not ( n2146 , n1447 ); 
or ( n2147 , n2145 , n2146 ); 
nand ( n2148 , n2142 , n1159 ); 
nand ( n2149 , n2147 , n2148 ); 
not ( n2150 , n2149 ); 
or ( n2151 , n2140 , n2150 ); 
nand ( n2152 , n2151 , n1175 ); 
nor ( n2153 , n2139 , n2152 ); 
not ( n2154 , n1321 ); 
not ( n2155 , n2144 ); 
not ( n2156 , n2155 ); 
or ( n2157 , n2154 , n2156 ); 
nand ( n2158 , n2157 , n67 ); 
or ( n2159 , n2153 , n2158 ); 
nand ( n2160 , n74 , n862 ); 
or ( n2161 , n67 , n2160 ); 
nand ( n2162 , n2159 , n2161 ); 
not ( n2163 , n1028 ); 
nand ( n2164 , n2163 , n1179 ); 
not ( n2165 , n860 ); 
not ( n2166 , n925 ); 
nor ( n2167 , n2166 , n890 ); 
xor ( n2168 , n2167 , n1371 ); 
nand ( n2169 , n2165 , n2168 ); 
and ( n2170 , n2164 , n2169 ); 
not ( n2171 , n959 ); 
nor ( n2172 , n992 , n1029 ); 
not ( n2173 , n2172 ); 
nand ( n2174 , n2173 , n1412 ); 
not ( n2175 , n1412 ); 
nand ( n2176 , n2172 , n2175 ); 
nand ( n2177 , n2171 , n2174 , n2176 ); 
not ( n2178 , n2177 ); 
nand ( n2179 , n2163 , n856 ); 
not ( n2180 , n2179 ); 
nor ( n2181 , n2178 , n2180 ); 
and ( n2182 , n2170 , n2181 ); 
not ( n2183 , n777 ); 
nor ( n2184 , n2182 , n2183 ); 
not ( n2185 , n1440 ); 
not ( n2186 , n77 ); 
nor ( n2187 , n2186 , n2 ); 
nand ( n2188 , n2187 , n956 ); 
nand ( n2189 , n2188 , n2169 , n2179 , n2177 ); 
not ( n2190 , n2189 ); 
not ( n2191 , n1842 ); 
or ( n2192 , n2190 , n2191 ); 
nand ( n2193 , n2187 , n1159 ); 
nand ( n2194 , n2192 , n2193 ); 
not ( n2195 , n2194 ); 
or ( n2196 , n2185 , n2195 ); 
nand ( n2197 , n2196 , n1175 ); 
nor ( n2198 , n2184 , n2197 ); 
not ( n2199 , n1993 ); 
not ( n2200 , n2189 ); 
not ( n2201 , n2200 ); 
or ( n2202 , n2199 , n2201 ); 
nand ( n2203 , n2202 , n67 ); 
or ( n2204 , n2198 , n2203 ); 
nand ( n2205 , n78 , n862 ); 
or ( n2206 , n67 , n2205 ); 
nand ( n2207 , n2204 , n2206 ); 
not ( n2208 , n971 ); 
nand ( n2209 , n2208 , n1636 ); 
not ( n2210 , n860 ); 
not ( n2211 , n945 ); 
nand ( n2212 , n2211 , n872 ); 
nand ( n2213 , n2212 , n1376 ); 
not ( n2214 , n2212 ); 
nand ( n2215 , n2214 , n1375 ); 
nand ( n2216 , n2210 , n2213 , n2215 ); 
and ( n2217 , n2209 , n2216 ); 
nand ( n2218 , n2208 , n1522 ); 
not ( n2219 , n2218 ); 
not ( n2220 , n959 ); 
not ( n2221 , n973 ); 
nor ( n2222 , n2221 , n1051 ); 
or ( n2223 , n2222 , n1422 ); 
nand ( n2224 , n2222 , n1422 ); 
nand ( n2225 , n2220 , n2223 , n2224 ); 
not ( n2226 , n2225 ); 
nor ( n2227 , n2219 , n2226 ); 
and ( n2228 , n2217 , n2227 ); 
nor ( n2229 , n2228 , n2183 ); 
not ( n2230 , n1575 ); 
not ( n2231 , n87 ); 
nor ( n2232 , n2231 , n2 ); 
nand ( n2233 , n2232 , n1206 ); 
nand ( n2234 , n2233 , n2216 , n2218 , n2225 ); 
not ( n2235 , n2234 ); 
not ( n2236 , n1842 ); 
or ( n2237 , n2235 , n2236 ); 
nand ( n2238 , n2232 , n1159 ); 
nand ( n2239 , n2237 , n2238 ); 
not ( n2240 , n2239 ); 
or ( n2241 , n2230 , n2240 ); 
nand ( n2242 , n2241 , n1175 ); 
nor ( n2243 , n2229 , n2242 ); 
not ( n2244 , n1453 ); 
not ( n2245 , n2234 ); 
not ( n2246 , n2245 ); 
or ( n2247 , n2244 , n2246 ); 
nand ( n2248 , n2247 , n67 ); 
or ( n2249 , n2243 , n2248 ); 
nand ( n2250 , n88 , n862 ); 
or ( n2251 , n67 , n2250 ); 
nand ( n2252 , n2249 , n2251 ); 
buf ( n2253 , n813 ); 
not ( n2254 , n2253 ); 
not ( n2255 , n2254 ); 
not ( n2256 , n1180 ); 
and ( n2257 , n2255 , n2256 ); 
not ( n2258 , n860 ); 
not ( n2259 , n936 ); 
nand ( n2260 , n2259 , n877 ); 
xor ( n2261 , n2260 , n1492 ); 
nand ( n2262 , n2258 , n2261 ); 
not ( n2263 , n2262 ); 
nor ( n2264 , n2257 , n2263 ); 
nand ( n2265 , n2253 , n856 ); 
not ( n2266 , n2265 ); 
not ( n2267 , n959 ); 
not ( n2268 , n981 ); 
nor ( n2269 , n2268 , n1042 ); 
buf ( n2270 , n1550 ); 
or ( n2271 , n2269 , n2270 ); 
nand ( n2272 , n2269 , n2270 ); 
nand ( n2273 , n2267 , n2271 , n2272 ); 
not ( n2274 , n2273 ); 
nor ( n2275 , n2266 , n2274 ); 
and ( n2276 , n2264 , n2275 ); 
nor ( n2277 , n2276 , n2183 ); 
not ( n2278 , n1575 ); 
not ( n2279 , n93 ); 
nor ( n2280 , n2279 , n2 ); 
nand ( n2281 , n2280 , n956 ); 
nand ( n2282 , n2281 , n2262 , n2265 , n2273 ); 
not ( n2283 , n2282 ); 
not ( n2284 , n1842 ); 
or ( n2285 , n2283 , n2284 ); 
nand ( n2286 , n2280 , n1159 ); 
nand ( n2287 , n2285 , n2286 ); 
not ( n2288 , n2287 ); 
or ( n2289 , n2278 , n2288 ); 
nand ( n2290 , n2289 , n1994 ); 
nor ( n2291 , n2277 , n2290 ); 
not ( n2292 , n1993 ); 
not ( n2293 , n2282 ); 
not ( n2294 , n2293 ); 
or ( n2295 , n2292 , n2294 ); 
nand ( n2296 , n2295 , n67 ); 
or ( n2297 , n2291 , n2296 ); 
nand ( n2298 , n94 , n862 ); 
or ( n2299 , n67 , n2298 ); 
nand ( n2300 , n2297 , n2299 ); 
nand ( n2301 , n99 , n862 ); 
not ( n2302 , n2301 ); 
nand ( n2303 , n2302 , n1179 ); 
not ( n2304 , n860 ); 
not ( n2305 , n943 ); 
nand ( n2306 , n2305 , n869 ); 
not ( n2307 , n938 ); 
nand ( n2308 , n2306 , n2307 ); 
not ( n2309 , n2306 ); 
nand ( n2310 , n2309 , n938 ); 
nand ( n2311 , n2304 , n2308 , n2310 ); 
buf ( n2312 , n942 ); 
nand ( n2313 , n2312 , n1601 ); 
not ( n2314 , n959 ); 
not ( n2315 , n968 ); 
nor ( n2316 , n2315 , n1048 ); 
xor ( n2317 , n2316 , n1044 ); 
nand ( n2318 , n2314 , n2317 ); 
nand ( n2319 , n2303 , n2311 , n2313 , n2318 ); 
not ( n2320 , n2319 ); 
not ( n2321 , n1626 ); 
or ( n2322 , n2320 , n2321 ); 
not ( n2323 , n2301 ); 
nand ( n2324 , n2323 , n1159 ); 
nand ( n2325 , n2322 , n2324 ); 
and ( n2326 , n2183 , n2325 ); 
not ( n2327 , n2312 ); 
not ( n2328 , n1179 ); 
or ( n2329 , n2327 , n2328 ); 
nand ( n2330 , n2329 , n2311 ); 
not ( n2331 , n2330 ); 
and ( n2332 , n2331 , n2313 , n2318 ); 
nor ( n2333 , n2332 , n1575 ); 
not ( n2334 , n1890 ); 
nor ( n2335 , n2326 , n2333 , n2334 ); 
not ( n2336 , n1321 ); 
not ( n2337 , n2319 ); 
not ( n2338 , n2337 ); 
or ( n2339 , n2336 , n2338 ); 
nand ( n2340 , n2339 , n67 ); 
or ( n2341 , n2335 , n2340 ); 
nand ( n2342 , n100 , n862 ); 
or ( n2343 , n67 , n2342 ); 
nand ( n2344 , n2341 , n2343 ); 
nand ( n2345 , n113 , n862 ); 
not ( n2346 , n2345 ); 
nor ( n2347 , n2346 , n776 ); 
and ( n2348 , n67 , n1192 ); 
not ( n2349 , n114 ); 
nor ( n2350 , n2349 , n2 ); 
not ( n2351 , n846 ); 
and ( n2352 , n2351 , n708 ); 
not ( n2353 , n558 ); 
nor ( n2354 , n2353 , n671 ); 
nand ( n2355 , n704 , n713 , n2354 , n494 ); 
nor ( n2356 , n2355 , n720 , n731 ); 
and ( n2357 , n707 , n2356 ); 
or ( n2358 , n707 , n2356 ); 
nand ( n2359 , n2358 , n846 ); 
nor ( n2360 , n2357 , n2359 ); 
nor ( n2361 , n2352 , n2360 ); 
not ( n2362 , n2361 ); 
and ( n2363 , n832 , n1167 ); 
nand ( n2364 , n741 , n769 ); 
nor ( n2365 , n2006 , n1958 ); 
and ( n2366 , n2365 , n804 , n800 ); 
and ( n2367 , n2366 , n611 , n664 , n817 ); 
and ( n2368 , n630 , n816 ); 
not ( n2369 , n1212 ); 
nor ( n2370 , n794 , n802 , n2369 ); 
nand ( n2371 , n2367 , n2368 , n1285 , n2370 ); 
nor ( n2372 , n2364 , n2371 ); 
not ( n2373 , n1508 ); 
nor ( n2374 , n2373 , n1081 ); 
and ( n2375 , n1510 , n340 ); 
not ( n2376 , n1855 ); 
and ( n2377 , n2375 , n2376 , n849 ); 
nand ( n2378 , n2363 , n2372 , n2374 , n2377 ); 
nand ( n2379 , n724 , n2378 ); 
not ( n2380 , n2379 ); 
nand ( n2381 , n2362 , n2380 ); 
not ( n2382 , n2381 ); 
not ( n2383 , n2382 ); 
nand ( n2384 , n2361 , n2379 ); 
nand ( n2385 , n2383 , n2384 ); 
not ( n2386 , n2351 ); 
or ( n2387 , n2386 , n711 ); 
not ( n2388 , n711 ); 
and ( n2389 , n704 , n707 , n838 , n756 ); 
not ( n2390 , n2389 ); 
or ( n2391 , n2388 , n2390 ); 
not ( n2392 , n711 ); 
not ( n2393 , n2389 ); 
and ( n2394 , n2392 , n2393 ); 
nor ( n2395 , n2394 , n2351 ); 
nand ( n2396 , n2391 , n2395 ); 
nand ( n2397 , n2387 , n2396 ); 
and ( n2398 , n2381 , n2397 ); 
not ( n2399 , n2381 ); 
not ( n2400 , n2397 ); 
and ( n2401 , n2399 , n2400 ); 
nor ( n2402 , n2398 , n2401 ); 
nand ( n2403 , n2350 , n2385 , n2402 ); 
not ( n2404 , n2402 ); 
nand ( n2405 , n2385 , n871 , n2404 ); 
and ( n2406 , n2403 , n2405 ); 
not ( n2407 , n2402 ); 
nor ( n2408 , n2407 , n2385 , n970 ); 
not ( n2409 , n2404 ); 
nor ( n2410 , n2160 , n2205 , n2298 , n2342 ); 
and ( n2411 , n2410 , n1901 , n1955 ); 
xor ( n2412 , n2411 , n2250 ); 
nor ( n2413 , n2409 , n2412 , n2385 ); 
nor ( n2414 , n2408 , n2413 ); 
nand ( n2415 , n776 , n2406 , n2414 ); 
nand ( n2416 , n2348 , n2415 ); 
or ( n2417 , n2347 , n2416 ); 
or ( n2418 , n2345 , n2348 ); 
nand ( n2419 , n2417 , n2418 ); 
or ( n2420 , n1339 , n849 ); 
nand ( n2421 , n206 , n862 ); 
not ( n2422 , n116 ); 
not ( n2423 , n862 ); 
or ( n2424 , n2422 , n2423 ); 
nand ( n2425 , n2424 , n1519 ); 
not ( n2426 , n2 ); 
nand ( n2427 , n2426 , n126 ); 
not ( n2428 , n2 ); 
nand ( n2429 , n2428 , n117 ); 
not ( n2430 , n2429 ); 
or ( n2431 , n2425 , n2427 , n2430 ); 
and ( n2432 , n118 , n862 ); 
nor ( n2433 , n2432 , n2055 , n1836 ); 
nor ( n2434 , n1722 , n1205 , n1442 , n1613 ); 
nand ( n2435 , n2433 , n2434 ); 
and ( n2436 , n1519 , n2435 ); 
and ( n2437 , n123 , n862 ); 
nor ( n2438 , n124 , n125 ); 
nor ( n2439 , n2 , n2438 ); 
nor ( n2440 , n2437 , n2439 ); 
and ( n2441 , n120 , n862 ); 
and ( n2442 , n119 , n862 ); 
nor ( n2443 , n2441 , n2442 ); 
and ( n2444 , n122 , n862 ); 
and ( n2445 , n121 , n862 ); 
nor ( n2446 , n2444 , n2445 ); 
and ( n2447 , n2440 , n2443 , n2446 ); 
nor ( n2448 , n2447 , n2427 ); 
nor ( n2449 , n2436 , n2448 ); 
and ( n2450 , n150 , n862 ); 
nor ( n2451 , n2450 , n1519 , n2429 ); 
not ( n2452 , n2430 ); 
nand ( n2453 , n135 , n136 ); 
nor ( n2454 , n2453 , n2 ); 
not ( n2455 , n2 ); 
nand ( n2456 , n2455 , n137 ); 
not ( n2457 , n2456 ); 
not ( n2458 , n138 ); 
nand ( n2459 , n139 , n140 , n141 ); 
nor ( n2460 , n2458 , n2459 , n2 ); 
nand ( n2461 , n2454 , n2457 , n2460 ); 
nand ( n2462 , n2452 , n2461 ); 
nand ( n2463 , n2449 , n2451 , n2427 , n2462 ); 
and ( n2464 , n2431 , n2463 ); 
or ( n2465 , n2421 , n2464 ); 
xor ( n2466 , n207 , n2421 ); 
not ( n2467 , n2 ); 
nand ( n2468 , n2467 , n115 ); 
not ( n2469 , n2468 ); 
nand ( n2470 , n2469 , n183 ); 
not ( n2471 , n183 ); 
nand ( n2472 , n2471 , n2468 ); 
not ( n2473 , n176 ); 
not ( n2474 , n2 ); 
nand ( n2475 , n2474 , n175 ); 
nand ( n2476 , n2473 , n2475 ); 
and ( n2477 , n2472 , n2476 ); 
not ( n2478 , n2477 ); 
not ( n2479 , n182 ); 
nor ( n2480 , n2479 , n2 ); 
nor ( n2481 , n181 , n2480 ); 
not ( n2482 , n2481 ); 
not ( n2483 , n177 ); 
not ( n2484 , n2 ); 
nand ( n2485 , n2484 , n178 ); 
nand ( n2486 , n2483 , n2485 ); 
nand ( n2487 , n2482 , n2486 ); 
nor ( n2488 , n2478 , n2487 ); 
not ( n2489 , n168 ); 
nor ( n2490 , n2489 , n2 ); 
or ( n2491 , n167 , n2490 ); 
not ( n2492 , n180 ); 
nor ( n2493 , n2492 , n2 ); 
or ( n2494 , n179 , n2493 ); 
and ( n2495 , n2491 , n2494 ); 
not ( n2496 , n2495 ); 
not ( n2497 , n170 ); 
nor ( n2498 , n2497 , n2 ); 
nor ( n2499 , n169 , n2498 ); 
not ( n2500 , n174 ); 
nor ( n2501 , n2500 , n2 ); 
nand ( n2502 , n173 , n2501 ); 
or ( n2503 , n2499 , n2502 ); 
nand ( n2504 , n169 , n2498 ); 
nand ( n2505 , n2503 , n2504 ); 
not ( n2506 , n2505 ); 
or ( n2507 , n2496 , n2506 ); 
not ( n2508 , n167 ); 
not ( n2509 , n2490 ); 
nor ( n2510 , n2508 , n2509 ); 
and ( n2511 , n2494 , n2510 ); 
nand ( n2512 , n179 , n2493 ); 
not ( n2513 , n2512 ); 
nor ( n2514 , n2511 , n2513 ); 
nand ( n2515 , n2507 , n2514 ); 
and ( n2516 , n2488 , n2515 ); 
nand ( n2517 , n181 , n2480 ); 
not ( n2518 , n2517 ); 
and ( n2519 , n2486 , n2518 ); 
not ( n2520 , n177 ); 
nor ( n2521 , n2520 , n2485 ); 
nor ( n2522 , n2519 , n2521 ); 
not ( n2523 , n2522 ); 
and ( n2524 , n2477 , n2523 ); 
nor ( n2525 , n2516 , n2524 ); 
nand ( n2526 , n2470 , n2525 ); 
not ( n2527 , n2472 ); 
not ( n2528 , n2475 ); 
nand ( n2529 , n2528 , n176 ); 
not ( n2530 , n2529 ); 
not ( n2531 , n2530 ); 
or ( n2532 , n2527 , n2531 ); 
not ( n2533 , n2495 ); 
nor ( n2534 , n173 , n2501 ); 
or ( n2535 , n2499 , n2534 ); 
nor ( n2536 , n2533 , n2535 ); 
not ( n2537 , n172 ); 
nor ( n2538 , n2537 , n2 ); 
or ( n2539 , n171 , n2538 ); 
not ( n2540 , n160 ); 
nor ( n2541 , n2540 , n2 ); 
nand ( n2542 , n159 , n2541 ); 
not ( n2543 , n2542 ); 
and ( n2544 , n2539 , n2543 ); 
nand ( n2545 , n171 , n2538 ); 
not ( n2546 , n2545 ); 
nor ( n2547 , n2544 , n2546 ); 
not ( n2548 , n2539 ); 
nor ( n2549 , n159 , n2541 ); 
nor ( n2550 , n2548 , n2549 ); 
not ( n2551 , n161 ); 
not ( n2552 , n2 ); 
nand ( n2553 , n2552 , n162 ); 
nand ( n2554 , n2551 , n2553 ); 
not ( n2555 , n164 ); 
nor ( n2556 , n2555 , n2 ); 
nand ( n2557 , n163 , n2556 ); 
not ( n2558 , n2557 ); 
and ( n2559 , n2554 , n2558 ); 
not ( n2560 , n2553 ); 
nand ( n2561 , n161 , n2560 ); 
not ( n2562 , n2561 ); 
nor ( n2563 , n2559 , n2562 ); 
not ( n2564 , n166 ); 
nor ( n2565 , n2564 , n2 ); 
nor ( n2566 , n165 , n2565 ); 
not ( n2567 , n156 ); 
nor ( n2568 , n2567 , n2 ); 
nand ( n2569 , n155 , n2568 ); 
or ( n2570 , n2566 , n2569 ); 
nand ( n2571 , n165 , n2565 ); 
nand ( n2572 , n2570 , n2571 ); 
not ( n2573 , n2572 ); 
not ( n2574 , n2573 ); 
not ( n2575 , n155 ); 
not ( n2576 , n2568 ); 
nand ( n2577 , n2575 , n2576 ); 
not ( n2578 , n2577 ); 
nor ( n2579 , n2578 , n2566 ); 
not ( n2580 , n152 ); 
nor ( n2581 , n2580 , n2 ); 
nor ( n2582 , n151 , n2581 ); 
not ( n2583 , n2582 ); 
not ( n2584 , n157 ); 
not ( n2585 , n158 ); 
nor ( n2586 , n2585 , n2 ); 
not ( n2587 , n2586 ); 
nand ( n2588 , n2584 , n2587 ); 
and ( n2589 , n2583 , n2588 ); 
not ( n2590 , n2589 ); 
not ( n2591 , n200 ); 
not ( n2592 , n201 ); 
nor ( n2593 , n2592 , n2 ); 
not ( n2594 , n2593 ); 
nand ( n2595 , n2591 , n2594 ); 
not ( n2596 , n2595 ); 
not ( n2597 , n203 ); 
nor ( n2598 , n2597 , n2 ); 
nand ( n2599 , n202 , n2598 ); 
not ( n2600 , n2599 ); 
not ( n2601 , n2600 ); 
or ( n2602 , n2596 , n2601 ); 
nand ( n2603 , n200 , n2593 ); 
nand ( n2604 , n2602 , n2603 ); 
not ( n2605 , n154 ); 
nor ( n2606 , n2605 , n2 ); 
nor ( n2607 , n153 , n2606 ); 
not ( n2608 , n199 ); 
nor ( n2609 , n2608 , n2 ); 
nor ( n2610 , n198 , n2609 ); 
nor ( n2611 , n2607 , n2610 ); 
and ( n2612 , n2604 , n2611 ); 
nand ( n2613 , n153 , n2606 ); 
nand ( n2614 , n198 , n2609 ); 
nand ( n2615 , n2613 , n2614 ); 
not ( n2616 , n2615 ); 
nand ( n2617 , n2613 , n2607 ); 
not ( n2618 , n2617 ); 
nor ( n2619 , n2616 , n2618 ); 
nor ( n2620 , n2612 , n2619 ); 
not ( n2621 , n205 ); 
nor ( n2622 , n2621 , n2 ); 
nor ( n2623 , n204 , n2622 ); 
not ( n2624 , n2 ); 
nand ( n2625 , n2624 , n191 ); 
not ( n2626 , n2625 ); 
nand ( n2627 , n190 , n2626 ); 
or ( n2628 , n2623 , n2627 ); 
nand ( n2629 , n204 , n2622 ); 
nand ( n2630 , n2628 , n2629 ); 
not ( n2631 , n2630 ); 
not ( n2632 , n190 ); 
nand ( n2633 , n2632 , n2625 ); 
not ( n2634 , n2633 ); 
nor ( n2635 , n2634 , n2623 ); 
not ( n2636 , n192 ); 
not ( n2637 , n2 ); 
nand ( n2638 , n2637 , n193 ); 
nand ( n2639 , n2636 , n2638 ); 
not ( n2640 , n2639 ); 
not ( n2641 , n195 ); 
nor ( n2642 , n2641 , n2 ); 
nand ( n2643 , n194 , n2642 ); 
not ( n2644 , n2643 ); 
not ( n2645 , n2644 ); 
or ( n2646 , n2640 , n2645 ); 
not ( n2647 , n2638 ); 
nand ( n2648 , n192 , n2647 ); 
nand ( n2649 , n2646 , n2648 ); 
nand ( n2650 , n2635 , n2649 ); 
not ( n2651 , n197 ); 
nor ( n2652 , n2651 , n2 ); 
nor ( n2653 , n196 , n2652 ); 
not ( n2654 , n185 ); 
nor ( n2655 , n2654 , n2 ); 
nand ( n2656 , n184 , n2655 ); 
or ( n2657 , n2653 , n2656 ); 
nand ( n2658 , n196 , n2652 ); 
nand ( n2659 , n2657 , n2658 ); 
not ( n2660 , n2659 ); 
not ( n2661 , n2660 ); 
not ( n2662 , n187 ); 
nor ( n2663 , n2662 , n2 ); 
and ( n2664 , n186 , n2663 ); 
not ( n2665 , n2664 ); 
not ( n2666 , n2665 ); 
not ( n2667 , n2 ); 
nand ( n2668 , n2667 , n188 ); 
not ( n2669 , n2668 ); 
not ( n2670 , n186 ); 
not ( n2671 , n2663 ); 
nand ( n2672 , n2670 , n2671 ); 
nand ( n2673 , n2669 , n189 , n2672 ); 
not ( n2674 , n2673 ); 
or ( n2675 , n2666 , n2674 ); 
not ( n2676 , n184 ); 
not ( n2677 , n2655 ); 
nand ( n2678 , n2676 , n2677 ); 
not ( n2679 , n2678 ); 
nor ( n2680 , n2679 , n2653 ); 
nand ( n2681 , n2675 , n2680 ); 
not ( n2682 , n2681 ); 
or ( n2683 , n2661 , n2682 ); 
not ( n2684 , n194 ); 
not ( n2685 , n2642 ); 
nand ( n2686 , n2684 , n2685 ); 
and ( n2687 , n2639 , n2686 ); 
and ( n2688 , n2687 , n2635 ); 
nand ( n2689 , n2683 , n2688 ); 
nand ( n2690 , n2631 , n2650 , n2689 ); 
not ( n2691 , n202 ); 
not ( n2692 , n2598 ); 
nand ( n2693 , n2691 , n2692 ); 
and ( n2694 , n2595 , n2693 ); 
nand ( n2695 , n2690 , n2611 , n2694 ); 
nand ( n2696 , n2620 , n2695 ); 
not ( n2697 , n2696 ); 
or ( n2698 , n2590 , n2697 ); 
nand ( n2699 , n151 , n2581 ); 
not ( n2700 , n2699 ); 
and ( n2701 , n2588 , n2700 ); 
nand ( n2702 , n157 , n2586 ); 
not ( n2703 , n2702 ); 
nor ( n2704 , n2701 , n2703 ); 
nand ( n2705 , n2698 , n2704 ); 
nand ( n2706 , n2579 , n2705 ); 
not ( n2707 , n2706 ); 
or ( n2708 , n2574 , n2707 ); 
or ( n2709 , n163 , n2556 ); 
and ( n2710 , n2554 , n2709 ); 
nand ( n2711 , n2708 , n2710 ); 
nand ( n2712 , n2563 , n2711 ); 
nand ( n2713 , n2550 , n2712 ); 
nand ( n2714 , n2547 , n2713 ); 
nand ( n2715 , n2536 , n2488 , n2714 ); 
nand ( n2716 , n2532 , n2715 ); 
nor ( n2717 , n2526 , n2716 ); 
or ( n2718 , n2466 , n2717 ); 
nand ( n2719 , n2466 , n2717 ); 
nand ( n2720 , n2718 , n2464 , n2719 ); 
nand ( n2721 , n2465 , n2720 ); 
nand ( n2722 , n1339 , n2721 ); 
nand ( n2723 , n2420 , n2722 ); 
or ( n2724 , n1339 , n832 ); 
or ( n2725 , n2468 , n2464 ); 
not ( n2726 , n2464 ); 
nor ( n2727 , n2582 , n2607 ); 
not ( n2728 , n2549 ); 
nand ( n2729 , n2728 , n2554 ); 
not ( n2730 , n2566 ); 
nand ( n2731 , n2730 , n2709 ); 
nor ( n2732 , n2729 , n2731 ); 
nand ( n2733 , n2577 , n2588 ); 
not ( n2734 , n2733 ); 
nand ( n2735 , n2599 , n2629 ); 
not ( n2736 , n2595 ); 
nor ( n2737 , n2736 , n2610 ); 
nor ( n2738 , n2600 , n2693 ); 
not ( n2739 , n2738 ); 
nand ( n2740 , n2735 , n2737 , n2739 ); 
or ( n2741 , n2610 , n2603 ); 
nand ( n2742 , n2741 , n2614 ); 
not ( n2743 , n2742 ); 
and ( n2744 , n2633 , n2639 ); 
not ( n2745 , n2686 ); 
or ( n2746 , n2745 , n2658 ); 
nand ( n2747 , n2746 , n2643 ); 
nand ( n2748 , n2744 , n2747 ); 
or ( n2749 , n2634 , n2648 ); 
nand ( n2750 , n2749 , n2627 ); 
not ( n2751 , n2750 ); 
nand ( n2752 , n2678 , n2664 ); 
nand ( n2753 , n2656 , n2752 ); 
nor ( n2754 , n2679 , n2673 ); 
or ( n2755 , n2753 , n2754 ); 
nor ( n2756 , n2745 , n2653 ); 
nand ( n2757 , n2755 , n2744 , n2756 ); 
nand ( n2758 , n2748 , n2751 , n2757 ); 
not ( n2759 , n2623 ); 
and ( n2760 , n2693 , n2759 ); 
nand ( n2761 , n2758 , n2737 , n2760 ); 
nand ( n2762 , n2740 , n2743 , n2761 ); 
nand ( n2763 , n2727 , n2732 , n2734 , n2762 ); 
not ( n2764 , n2491 ); 
nor ( n2765 , n2764 , n2499 ); 
not ( n2766 , n2539 ); 
nor ( n2767 , n2766 , n2534 ); 
nand ( n2768 , n2765 , n2767 ); 
not ( n2769 , n2481 ); 
nand ( n2770 , n2769 , n2494 ); 
not ( n2771 , n2770 ); 
and ( n2772 , n2476 , n2486 ); 
nand ( n2773 , n2771 , n2772 ); 
nor ( n2774 , n2763 , n2768 , n2773 ); 
or ( n2775 , n2481 , n2512 ); 
nand ( n2776 , n2775 , n2517 ); 
and ( n2777 , n2772 , n2776 ); 
and ( n2778 , n2476 , n2521 ); 
nor ( n2779 , n2777 , n2778 ); 
not ( n2780 , n2779 ); 
not ( n2781 , n2768 ); 
or ( n2782 , n2549 , n2561 ); 
nand ( n2783 , n2782 , n2542 ); 
not ( n2784 , n2783 ); 
not ( n2785 , n2729 ); 
not ( n2786 , n2709 ); 
or ( n2787 , n2786 , n2571 ); 
nand ( n2788 , n2787 , n2557 ); 
nand ( n2789 , n2785 , n2788 ); 
not ( n2790 , n2699 ); 
not ( n2791 , n2582 ); 
or ( n2792 , n2790 , n2791 ); 
nand ( n2793 , n2699 , n2613 ); 
nand ( n2794 , n2792 , n2793 ); 
or ( n2795 , n2733 , n2794 ); 
or ( n2796 , n2578 , n2702 ); 
nand ( n2797 , n2796 , n2569 ); 
not ( n2798 , n2797 ); 
nand ( n2799 , n2795 , n2798 ); 
nand ( n2800 , n2732 , n2799 ); 
nand ( n2801 , n2784 , n2789 , n2800 ); 
and ( n2802 , n2781 , n2801 ); 
not ( n2803 , n2765 ); 
or ( n2804 , n2534 , n2545 ); 
nand ( n2805 , n2804 , n2502 ); 
not ( n2806 , n2805 ); 
or ( n2807 , n2803 , n2806 ); 
not ( n2808 , n2504 ); 
and ( n2809 , n2491 , n2808 ); 
nor ( n2810 , n2809 , n2510 ); 
nand ( n2811 , n2807 , n2810 ); 
nor ( n2812 , n2802 , n2811 ); 
or ( n2813 , n2773 , n2812 ); 
nand ( n2814 , n2813 , n2529 ); 
nor ( n2815 , n2780 , n2814 ); 
not ( n2816 , n2815 ); 
or ( n2817 , n2774 , n2816 ); 
nand ( n2818 , n2472 , n2470 ); 
nand ( n2819 , n2817 , n2818 ); 
or ( n2820 , n2726 , n2819 ); 
not ( n2821 , n2818 ); 
not ( n2822 , n2774 ); 
nand ( n2823 , n2821 , n2822 , n2464 , n2815 ); 
nand ( n2824 , n2725 , n2820 , n2823 ); 
nand ( n2825 , n1339 , n2824 ); 
nand ( n2826 , n2724 , n2825 ); 
not ( n2827 , n832 ); 
not ( n2828 , n1339 ); 
or ( n2829 , n2475 , n2464 ); 
and ( n2830 , n2694 , n2635 ); 
not ( n2831 , n2681 ); 
and ( n2832 , n2830 , n2687 , n2831 ); 
nor ( n2833 , n2832 , n2604 ); 
not ( n2834 , n2649 ); 
nand ( n2835 , n2687 , n2659 ); 
nand ( n2836 , n2834 , n2835 ); 
and ( n2837 , n2830 , n2836 ); 
and ( n2838 , n2694 , n2630 ); 
nor ( n2839 , n2837 , n2838 ); 
and ( n2840 , n2833 , n2839 ); 
not ( n2841 , n2487 ); 
nand ( n2842 , n2841 , n2495 ); 
not ( n2843 , n2842 ); 
not ( n2844 , n2550 ); 
nor ( n2845 , n2844 , n2535 ); 
nand ( n2846 , n2843 , n2589 , n2611 , n2845 ); 
nand ( n2847 , n2710 , n2579 ); 
nor ( n2848 , n2840 , n2846 , n2847 ); 
or ( n2849 , n2487 , n2514 ); 
nand ( n2850 , n2710 , n2572 ); 
not ( n2851 , n2847 ); 
nand ( n2852 , n2617 , n2615 , n2589 ); 
nand ( n2853 , n2704 , n2852 ); 
nand ( n2854 , n2851 , n2853 ); 
nand ( n2855 , n2563 , n2850 , n2854 ); 
and ( n2856 , n2845 , n2855 ); 
nor ( n2857 , n2535 , n2547 ); 
nor ( n2858 , n2856 , n2505 , n2857 ); 
or ( n2859 , n2842 , n2858 ); 
nand ( n2860 , n2849 , n2859 , n2522 ); 
or ( n2861 , n2848 , n2860 ); 
nand ( n2862 , n2476 , n2529 ); 
nand ( n2863 , n2861 , n2862 ); 
or ( n2864 , n2726 , n2863 ); 
not ( n2865 , n2848 ); 
not ( n2866 , n2860 ); 
not ( n2867 , n2862 ); 
nand ( n2868 , n2865 , n2464 , n2866 , n2867 ); 
nand ( n2869 , n2829 , n2864 , n2868 ); 
not ( n2870 , n2869 ); 
or ( n2871 , n2828 , n2870 ); 
or ( n2872 , n1339 , n770 ); 
nand ( n2873 , n2871 , n2872 ); 
not ( n2874 , n1339 ); 
or ( n2875 , n2485 , n2464 ); 
and ( n2876 , n2744 , n2760 ); 
nand ( n2877 , n2876 , n2756 , n2754 ); 
and ( n2878 , n2756 , n2753 ); 
or ( n2879 , n2747 , n2878 ); 
nand ( n2880 , n2879 , n2876 ); 
and ( n2881 , n2750 , n2760 ); 
not ( n2882 , n2735 ); 
nor ( n2883 , n2882 , n2738 ); 
nor ( n2884 , n2881 , n2883 ); 
and ( n2885 , n2877 , n2880 , n2884 ); 
not ( n2886 , n2770 ); 
nand ( n2887 , n2886 , n2765 ); 
nor ( n2888 , n2885 , n2887 ); 
nand ( n2889 , n2888 , n2727 , n2737 ); 
not ( n2890 , n2731 ); 
nand ( n2891 , n2890 , n2734 ); 
nand ( n2892 , n2785 , n2767 ); 
nor ( n2893 , n2889 , n2891 , n2892 ); 
or ( n2894 , n2770 , n2810 ); 
not ( n2895 , n2892 ); 
and ( n2896 , n2727 , n2742 ); 
not ( n2897 , n2794 ); 
nor ( n2898 , n2896 , n2897 ); 
or ( n2899 , n2891 , n2898 ); 
or ( n2900 , n2731 , n2798 ); 
not ( n2901 , n2788 ); 
nand ( n2902 , n2899 , n2900 , n2901 ); 
and ( n2903 , n2895 , n2902 ); 
and ( n2904 , n2767 , n2783 ); 
nor ( n2905 , n2903 , n2904 , n2805 ); 
or ( n2906 , n2887 , n2905 ); 
not ( n2907 , n2776 ); 
nand ( n2908 , n2894 , n2906 , n2907 ); 
or ( n2909 , n2893 , n2908 ); 
not ( n2910 , n2521 ); 
nand ( n2911 , n2910 , n2486 ); 
nand ( n2912 , n2909 , n2911 ); 
or ( n2913 , n2726 , n2912 ); 
not ( n2914 , n2911 ); 
not ( n2915 , n2908 ); 
not ( n2916 , n2893 ); 
nand ( n2917 , n2914 , n2464 , n2915 , n2916 ); 
nand ( n2918 , n2875 , n2913 , n2917 ); 
not ( n2919 , n2918 ); 
or ( n2920 , n2874 , n2919 ); 
or ( n2921 , n1339 , n741 ); 
nand ( n2922 , n2920 , n2921 ); 
patch p0 (.t_0(t_0), .g1(n555), .g2(n550), .g3(n545));
endmodule 

