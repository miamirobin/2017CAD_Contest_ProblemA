module patch (t_0, t_1, t_2, t_3, g1, g2, g3, g4, g5, g6, g7, g8);
input g1, g2, g3, g4, g5, g6, g7, g8;
output t_0, t_1, t_2, t_3;
wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237;

and ( w1 , g2 , g3 );
and ( w2 , w183 , w1 );
and ( w3 , w2 , g4 );
and ( w4 , w3 , w188 );
and ( w5 , w4 , w134 );
and ( w6 , g7 , w226 );
and ( w7 , w6 , g5 );
and ( w8 , w7 , g3 );
and ( w9 , w8 , g6 );
nor ( w10 , w5 , w9 );
and ( w11 , g7 , g6 );
not ( w12 , w8 );
and ( w13 , w11 , w12 );
and ( w14 , g6 , w226 );
and ( w15 , w148 , g3 );
nor ( w16 , w13 , w15 );
and ( w17 , w16 , g5 );
and ( w18 , w17 , g3 );
nor ( w19 , g6 , g5 );
nor ( w20 , g2 , g3 );
nor ( w21 , w20 , w1 );
and ( w22 , w19 , w39 );
and ( w23 , w22 , g4 );
not ( w24 , w23 );
and ( w25 , w10 , w24 );
nor ( w26 , w25 , g3 );
nor ( w27 , g7 , w26 );
nor ( w28 , w27 , g6 );
and ( w29 , w28 , w188 );
and ( w30 , w29 , g2 );
nor ( w31 , w30 , w23 );
nor ( w32 , w31 , g3 );
nor ( w33 , w18 , w32 );
nor ( w34 , w33 , g4 );
and ( w35 , w183 , g4 );
and ( w36 , w35 , w188 );
and ( w37 , w36 , g3 );
and ( w38 , w37 , g6 );
not ( w39 , w21 );
and ( w40 , w38 , w39 );
and ( w41 , w40 , g3 );
nor ( w42 , w41 , w32 );
not ( w43 , w34 );
and ( w44 , w43 , w42 );
nand ( t_0 , w10 , w44 );
and ( w45 , g3 , g7 );
and ( w46 , w45 , w134 );
nor ( w47 , g7 , g3 );
and ( w48 , w47 , g6 );
and ( w49 , w48 , w21 );
nor ( w50 , w49 , w5 );
and ( w51 , w21 , w228 );
nor ( w52 , w51 , g6 );
not ( w53 , w52 );
and ( w54 , w53 , g7 );
and ( w55 , w54 , w21 );
and ( w56 , w55 , w188 );
and ( w57 , w134 , w56 );
nor ( w58 , w57 , w5 );
and ( w59 , w14 , w228 );
nor ( w60 , w4 , w59 );
not ( w61 , w60 );
and ( w62 , w61 , g4 );
and ( w63 , w62 , w188 );
not ( w64 , w63 );
and ( w65 , w58 , w64 );
and ( w66 , w50 , w65 );
nor ( w67 , w66 , g4 );
not ( w68 , w67 );
and ( w69 , w68 , w65 );
not ( w70 , w69 );
and ( w71 , w70 , g5 );
nor ( w72 , w71 , w5 );
and ( w73 , w72 , w65 );
not ( w74 , w46 );
and ( w75 , w74 , w73 );
not ( w76 , w75 );
and ( w77 , w76 , w21 );
not ( w78 , w77 );
and ( w79 , w78 , w73 );
not ( w80 , w79 );
and ( w81 , w80 , g5 );
not ( w82 , w81 );
and ( w83 , w82 , w73 );
and ( w84 , w153 , g6 );
and ( w85 , w84 , g3 );
and ( w86 , w49 , w102 );
and ( w87 , w86 , g5 );
nor ( w88 , w85 , w87 );
not ( w89 , w88 );
and ( w90 , w89 , w21 );
and ( w91 , w90 , w102 );
and ( w92 , w91 , g5 );
not ( w93 , w92 );
and ( w94 , w83 , w93 );
and ( w95 , w94 , w134 );
nor ( w96 , w95 , g2 );
not ( w97 , w96 );
and ( w98 , w94 , w97 );
not ( w99 , w98 );
and ( w100 , w99 , g4 );
and ( w101 , w134 , w21 );
not ( w102 , g4 );
and ( w103 , w101 , w102 );
not ( w104 , w103 );
and ( w105 , w104 , w94 );
nor ( w106 , w105 , g3 );
and ( w107 , w106 , w188 );
nor ( w108 , w100 , w107 );
nor ( w109 , w108 , g3 );
not ( w110 , w109 );
and ( w111 , w110 , w94 );
nor ( w112 , w111 , g5 );
and ( t_1 , w94 , w237 );
nor ( w113 , g5 , g7 );
and ( w114 , w113 , g6 );
and ( w115 , w114 , g2 );
and ( w116 , w115 , w228 );
nor ( w117 , w116 , g7 );
and ( w118 , w117 , g2 );
and ( w119 , g2 , w134 );
nor ( w120 , w119 , w14 );
nor ( w121 , w120 , g3 );
not ( w122 , w121 );
and ( w123 , w118 , w122 );
not ( w124 , w113 );
and ( w125 , w124 , g6 );
nor ( w126 , w125 , g4 );
and ( w127 , w126 , w228 );
nor ( w128 , w127 , w121 );
nor ( w129 , g2 , g6 );
and ( w130 , w188 , g2 );
and ( w131 , w130 , g6 );
nor ( w132 , w131 , g3 );
and ( w133 , w226 , g3 );
not ( w134 , g6 );
and ( w135 , w133 , w134 );
nor ( w136 , w132 , w135 );
nor ( w137 , w129 , w136 );
and ( w138 , w137 , g4 );
nor ( w139 , w138 , w14 );
nor ( w140 , w139 , g3 );
nor ( w141 , w140 , w135 );
nor ( w142 , w121 , w14 );
nor ( w143 , w142 , g3 );
not ( w144 , w143 );
and ( w145 , w141 , w144 );
and ( w146 , w145 , g8 );
and ( w147 , w146 , w153 );
not ( w148 , w14 );
and ( w149 , w147 , w148 );
nor ( w150 , w149 , g3 );
nor ( w151 , w150 , w135 );
and ( w152 , w128 , w151 );
not ( w153 , g7 );
and ( w154 , w152 , w153 );
and ( w155 , w154 , g4 );
and ( w156 , w155 , w228 );
nor ( w157 , w156 , g2 );
and ( w158 , g6 , g2 );
nor ( w159 , w158 , g3 );
not ( w160 , w157 );
and ( w161 , w160 , w159 );
and ( w162 , w121 , w226 );
nor ( w163 , w162 , g3 );
not ( w164 , w158 );
and ( w165 , w164 , w163 );
and ( w166 , w165 , w188 );
and ( w167 , w166 , g7 );
and ( w168 , w154 , w228 );
nor ( w169 , w167 , w168 );
not ( w170 , w169 );
and ( w171 , w161 , w170 );
and ( w172 , w171 , w188 );
nor ( w173 , w123 , w172 );
nor ( w174 , w173 , g4 );
nor ( w175 , w174 , w172 );
nor ( w176 , w175 , w169 );
nor ( w177 , w1 , g5 );
not ( w178 , w20 );
and ( w179 , w178 , w177 );
nor ( w180 , w179 , g5 );
and ( w181 , g3 , w180 );
and ( w182 , w181 , g6 );
not ( w183 , g1 );
and ( w184 , w182 , w183 );
and ( w185 , w184 , g4 );
and ( w186 , w185 , w188 );
nor ( w187 , w176 , w186 );
not ( w188 , g5 );
and ( w189 , w188 , w187 );
and ( w190 , w135 , g7 );
and ( w191 , g6 , w21 );
nor ( w192 , w129 , w191 );
nor ( w193 , w192 , g2 );
and ( w194 , w193 , g6 );
nor ( w195 , w194 , w49 );
not ( w196 , w176 );
and ( w197 , w195 , w196 );
nor ( w198 , w197 , g7 );
and ( w199 , g6 , w20 );
nor ( w200 , w199 , w101 );
and ( w201 , w200 , w228 );
and ( w202 , w201 , g6 );
and ( w203 , w202 , g7 );
not ( w204 , w203 );
and ( w205 , w204 , w187 );
not ( w206 , w205 );
and ( w207 , w206 , g5 );
not ( w208 , w207 );
and ( w209 , w208 , w187 );
not ( w210 , w198 );
and ( w211 , w210 , w209 );
nor ( w212 , w211 , g4 );
not ( w213 , w212 );
and ( w214 , w213 , w187 );
not ( w215 , w214 );
and ( w216 , w215 , g5 );
not ( w217 , w216 );
and ( w218 , w217 , w187 );
not ( w219 , w190 );
and ( w220 , w219 , w218 );
not ( w221 , w220 );
and ( w222 , w221 , g5 );
not ( w223 , w222 );
and ( w224 , w223 , w187 );
and ( w225 , g6 , w224 );
not ( w226 , g2 );
and ( w227 , w226 , w224 );
not ( w228 , g3 );
and ( w229 , w228 , w224 );
nor ( w230 , w227 , w229 );
not ( w231 , w225 );
and ( w232 , w231 , w230 );
not ( w233 , w189 );
and ( w234 , w233 , w232 );
and ( w235 , w234 , g7 );
not ( w236 , w235 );
nand ( t_2 , w236 , w224 );
not ( w237 , w112 );
and ( t_3 , w94 , w237 );

endmodule
