module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 ); 
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 ; 
output g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 ; 

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 ; 
wire t_0 ; 
buf ( n1 , g0 ); 
buf ( n2 , g1 ); 
buf ( n3 , g2 ); 
buf ( n4 , g3 ); 
buf ( n5 , g4 ); 
buf ( n6 , g5 ); 
buf ( n7 , g6 ); 
buf ( n8 , g7 ); 
buf ( n9 , g8 ); 
buf ( n10 , g9 ); 
buf ( n11 , g10 ); 
buf ( n12 , g11 ); 
buf ( n13 , g12 ); 
buf ( n14 , g13 ); 
buf ( n15 , g14 ); 
buf ( n16 , g15 ); 
buf ( n17 , g16 ); 
buf ( n18 , g17 ); 
buf ( n19 , g18 ); 
buf ( n20 , g19 ); 
buf ( n21 , g20 ); 
buf ( n22 , g21 ); 
buf ( n23 , g22 ); 
buf ( n24 , g23 ); 
buf ( n25 , g24 ); 
buf ( n26 , g25 ); 
buf ( n27 , g26 ); 
buf ( n28 , g27 ); 
buf ( n29 , g28 ); 
buf ( n30 , g29 ); 
buf ( n31 , g30 ); 
buf ( n32 , g31 ); 
buf ( n33 , g32 ); 
buf ( n34 , g33 ); 
buf ( n35 , g34 ); 
buf ( n36 , g35 ); 
buf ( n37 , g36 ); 
buf ( n38 , g37 ); 
buf ( n39 , g38 ); 
buf ( n40 , g39 ); 
buf ( n41 , g40 ); 
buf ( n42 , g41 ); 
buf ( n43 , g42 ); 
buf ( n44 , g43 ); 
buf ( n45 , g44 ); 
buf ( n46 , g45 ); 
buf ( n47 , g46 ); 
buf ( n48 , g47 ); 
buf ( n49 , g48 ); 
buf ( n50 , g49 ); 
buf ( n51 , g50 ); 
buf ( n52 , g51 ); 
buf ( n53 , g52 ); 
buf ( n54 , g53 ); 
buf ( n55 , g54 ); 
buf ( n56 , g55 ); 
buf ( n57 , g56 ); 
buf ( n58 , g57 ); 
buf ( n59 , g58 ); 
buf ( n60 , g59 ); 
buf ( n61 , g60 ); 
buf ( n62 , g61 ); 
buf ( n63 , g62 ); 
buf ( n64 , g63 ); 
buf ( n65 , g64 ); 
buf ( n66 , g65 ); 
buf ( n67 , g66 ); 
buf ( n68 , g67 ); 
buf ( n69 , g68 ); 
buf ( n70 , g69 ); 
buf ( n71 , g70 ); 
buf ( n72 , g71 ); 
buf ( n73 , g72 ); 
buf ( n74 , g73 ); 
buf ( n75 , g74 ); 
buf ( n76 , g75 ); 
buf ( n77 , g76 ); 
buf ( n78 , g77 ); 
buf ( n79 , g78 ); 
buf ( n80 , g79 ); 
buf ( n81 , g80 ); 
buf ( n82 , g81 ); 
buf ( n83 , g82 ); 
buf ( n84 , g83 ); 
buf ( n85 , g84 ); 
buf ( n86 , g85 ); 
buf ( n87 , g86 ); 
buf ( n88 , g87 ); 
buf ( n89 , g88 ); 
buf ( n90 , g89 ); 
buf ( n91 , g90 ); 
buf ( n92 , g91 ); 
buf ( n93 , g92 ); 
buf ( n94 , g93 ); 
buf ( n95 , g94 ); 
buf ( n96 , g95 ); 
buf ( n97 , g96 ); 
buf ( n98 , g97 ); 
buf ( n99 , g98 ); 
buf ( n100 , g99 ); 
buf ( n101 , g100 ); 
buf ( n102 , g101 ); 
buf ( n103 , g102 ); 
buf ( n104 , g103 ); 
buf ( n105 , g104 ); 
buf ( n106 , g105 ); 
buf ( n107 , g106 ); 
buf ( n108 , g107 ); 
buf ( n109 , g108 ); 
buf ( n110 , g109 ); 
buf ( n111 , g110 ); 
buf ( n112 , g111 ); 
buf ( n113 , g112 ); 
buf ( n114 , g113 ); 
buf ( n115 , g114 ); 
buf ( n116 , g115 ); 
buf ( n117 , g116 ); 
buf ( n118 , g117 ); 
buf ( n119 , g118 ); 
buf ( n120 , g119 ); 
buf ( n121 , g120 ); 
buf ( n122 , g121 ); 
buf ( n123 , g122 ); 
buf ( n124 , g123 ); 
buf ( n125 , g124 ); 
buf ( n126 , g125 ); 
buf ( n127 , g126 ); 
buf ( n128 , g127 ); 
buf ( n129 , g128 ); 
buf ( n130 , g129 ); 
buf ( n131 , g130 ); 
buf ( n132 , g131 ); 
buf ( n133 , g132 ); 
buf ( n134 , g133 ); 
buf ( n135 , g134 ); 
buf ( n136 , g135 ); 
buf ( n137 , g136 ); 
buf ( n138 , g137 ); 
buf ( n139 , g138 ); 
buf ( n140 , g139 ); 
buf ( n141 , g140 ); 
buf ( n142 , g141 ); 
buf ( n143 , g142 ); 
buf ( n144 , g143 ); 
buf ( n145 , g144 ); 
buf ( n146 , g145 ); 
buf ( n147 , g146 ); 
buf ( n148 , g147 ); 
buf ( n149 , g148 ); 
buf ( n150 , g149 ); 
buf ( n151 , g150 ); 
buf ( n152 , g151 ); 
buf ( n153 , g152 ); 
buf ( n154 , g153 ); 
buf ( n155 , g154 ); 
buf ( n156 , g155 ); 
buf ( n157 , g156 ); 
buf ( n158 , g157 ); 
buf ( n159 , g158 ); 
buf ( n160 , g159 ); 
buf ( n161 , g160 ); 
buf ( n162 , g161 ); 
buf ( n163 , g162 ); 
buf ( n164 , g163 ); 
buf ( n165 , g164 ); 
buf ( n166 , g165 ); 
buf ( n167 , g166 ); 
buf ( n168 , g167 ); 
buf ( n169 , g168 ); 
buf ( n170 , g169 ); 
buf ( n171 , g170 ); 
buf ( n172 , g171 ); 
buf ( n173 , g172 ); 
buf ( n174 , g173 ); 
buf ( n175 , g174 ); 
buf ( n176 , g175 ); 
buf ( n177 , g176 ); 
buf ( n178 , g177 ); 
buf ( n179 , g178 ); 
buf ( n180 , g179 ); 
buf ( n181 , g180 ); 
buf ( n182 , g181 ); 
buf ( n183 , g182 ); 
buf ( n184 , g183 ); 
buf ( n185 , g184 ); 
buf ( n186 , g185 ); 
buf ( n187 , g186 ); 
buf ( n188 , g187 ); 
buf ( n189 , g188 ); 
buf ( n190 , g189 ); 
buf ( n191 , g190 ); 
buf ( n192 , g191 ); 
buf ( n193 , g192 ); 
buf ( n194 , g193 ); 
buf ( n195 , g194 ); 
buf ( n196 , g195 ); 
buf ( n197 , g196 ); 
buf ( n198 , g197 ); 
buf ( g198 , n199 ); 
buf ( g199 , n200 ); 
buf ( g200 , n201 ); 
buf ( g201 , n202 ); 
buf ( g202 , n203 ); 
buf ( g203 , n204 ); 
buf ( g204 , n205 ); 
buf ( g205 , n206 ); 
buf ( g206 , n207 ); 
buf ( g207 , n208 ); 
buf ( g208 , n209 ); 
buf ( g209 , n210 ); 
buf ( g210 , n211 ); 
buf ( g211 , n212 ); 
buf ( n199 , n1312 ); 
buf ( n200 , n1872 ); 
buf ( n201 , n1870 ); 
buf ( n202 , n1668 ); 
buf ( n203 , n1327 ); 
buf ( n204 , n865 ); 
buf ( n205 , n1871 ); 
buf ( n206 , n873 ); 
buf ( n207 , n873 ); 
buf ( n208 , n1502 ); 
buf ( n209 , n67 ); 
buf ( n210 , n70 ); 
buf ( n211 , n73 ); 
buf ( n212 , n78 ); 
not ( n216 , n120 ); 
nand ( n217 , n1 , n216 ); 
not ( n218 , n119 ); 
nand ( n219 , n218 , n1 ); 
not ( n220 , n219 ); 
and ( n221 , n217 , n3 ); 
not ( n222 , n217 ); 
not ( n223 , n3 ); 
and ( n224 , n222 , n223 ); 
nor ( n225 , n221 , n224 ); 
not ( n226 , n225 ); 
nor ( n227 , n220 , n226 ); 
or ( n228 , n217 , n227 ); 
nand ( n229 , n228 , n3 ); 
and ( n230 , n6 , n10 ); 
not ( n231 , n6 ); 
not ( n232 , n126 ); 
and ( n233 , n231 , n232 ); 
nor ( n234 , n230 , n233 ); 
not ( n235 , n234 ); 
not ( n236 , n235 ); 
not ( n237 , n6 ); 
not ( n238 , n166 ); 
not ( n239 , n238 ); 
or ( n240 , n237 , n239 ); 
nand ( n241 , n8 , n9 ); 
buf ( n242 , n241 ); 
nand ( n243 , n240 , n242 ); 
and ( n244 , n236 , n243 ); 
not ( n245 , n236 ); 
not ( n246 , n243 ); 
and ( n247 , n245 , n246 ); 
or ( n248 , n244 , n247 ); 
not ( n249 , n6 ); 
not ( n250 , n165 ); 
not ( n251 , n250 ); 
or ( n252 , n249 , n251 ); 
nand ( n253 , n8 , n9 ); 
buf ( n254 , n253 ); 
nand ( n255 , n252 , n254 ); 
not ( n256 , n255 ); 
not ( n257 , n256 ); 
and ( n258 , n6 , n12 ); 
not ( n259 , n6 ); 
not ( n260 , n125 ); 
and ( n261 , n259 , n260 ); 
nor ( n262 , n258 , n261 ); 
not ( n263 , n262 ); 
not ( n264 , n263 ); 
or ( n265 , n257 , n264 ); 
or ( n266 , n256 , n263 ); 
nand ( n267 , n265 , n266 ); 
and ( n268 , n248 , n267 ); 
not ( n269 , n6 ); 
not ( n270 , n167 ); 
not ( n271 , n270 ); 
or ( n272 , n269 , n271 ); 
nand ( n273 , n272 , n242 ); 
not ( n274 , n273 ); 
not ( n275 , n274 ); 
and ( n276 , n6 , n5 ); 
not ( n277 , n6 ); 
not ( n278 , n127 ); 
and ( n279 , n277 , n278 ); 
nor ( n280 , n276 , n279 ); 
not ( n281 , n280 ); 
not ( n282 , n281 ); 
or ( n283 , n275 , n282 ); 
nand ( n284 , n273 , n280 ); 
nand ( n285 , n283 , n284 ); 
not ( n286 , n254 ); 
not ( n287 , n286 ); 
and ( n288 , n6 , n16 ); 
not ( n289 , n6 ); 
not ( n290 , n123 ); 
and ( n291 , n289 , n290 ); 
nor ( n292 , n288 , n291 ); 
nand ( n293 , n287 , n292 ); 
not ( n294 , n287 ); 
not ( n295 , n292 ); 
and ( n296 , n294 , n295 ); 
not ( n297 , n6 ); 
not ( n298 , n164 ); 
not ( n299 , n298 ); 
or ( n300 , n297 , n299 ); 
nand ( n301 , n300 , n254 ); 
not ( n302 , n301 ); 
not ( n303 , n14 ); 
and ( n304 , n6 , n303 ); 
not ( n305 , n6 ); 
and ( n306 , n305 , n124 ); 
nor ( n307 , n304 , n306 ); 
not ( n308 , n307 ); 
not ( n309 , n308 ); 
and ( n310 , n302 , n309 ); 
and ( n311 , n301 , n308 ); 
nor ( n312 , n310 , n311 ); 
nor ( n313 , n296 , n312 ); 
and ( n314 , n268 , n285 , n293 , n313 ); 
not ( n315 , n314 ); 
and ( n316 , n6 , n181 ); 
not ( n317 , n6 ); 
and ( n318 , n317 , n42 ); 
or ( n319 , n316 , n318 ); 
not ( n320 , n319 ); 
and ( n321 , n6 , n40 ); 
not ( n322 , n6 ); 
not ( n323 , n142 ); 
and ( n324 , n322 , n323 ); 
nor ( n325 , n321 , n324 ); 
nand ( n326 , n320 , n325 ); 
not ( n327 , n325 ); 
nand ( n328 , n319 , n327 ); 
nand ( n329 , n326 , n328 ); 
not ( n330 , n43 ); 
and ( n331 , n6 , n330 ); 
not ( n332 , n6 ); 
and ( n333 , n332 , n141 ); 
nor ( n334 , n331 , n333 ); 
not ( n335 , n334 ); 
not ( n336 , n335 ); 
and ( n337 , n6 , n180 ); 
not ( n338 , n6 ); 
and ( n339 , n338 , n45 ); 
nor ( n340 , n337 , n339 ); 
not ( n341 , n340 ); 
and ( n342 , n336 , n341 ); 
and ( n343 , n340 , n335 ); 
nor ( n344 , n342 , n343 ); 
not ( n345 , n344 ); 
and ( n346 , n6 , n179 ); 
not ( n347 , n6 ); 
and ( n348 , n347 , n48 ); 
nor ( n349 , n346 , n348 ); 
not ( n350 , n349 ); 
and ( n351 , n6 , n46 ); 
not ( n352 , n6 ); 
not ( n353 , n140 ); 
and ( n354 , n352 , n353 ); 
nor ( n355 , n351 , n354 ); 
not ( n356 , n355 ); 
or ( n357 , n350 , n356 ); 
not ( n358 , n349 ); 
not ( n359 , n355 ); 
nand ( n360 , n358 , n359 ); 
nand ( n361 , n357 , n360 ); 
and ( n362 , n6 , n51 ); 
not ( n363 , n6 ); 
not ( n364 , n139 ); 
and ( n365 , n363 , n364 ); 
nor ( n366 , n362 , n365 ); 
not ( n367 , n366 ); 
not ( n368 , n6 ); 
not ( n369 , n178 ); 
or ( n370 , n368 , n369 ); 
not ( n371 , n6 ); 
nand ( n372 , n371 , n50 ); 
nand ( n373 , n370 , n372 ); 
not ( n374 , n373 ); 
and ( n375 , n367 , n374 ); 
not ( n376 , n367 ); 
and ( n377 , n376 , n373 ); 
nor ( n378 , n375 , n377 ); 
and ( n379 , n329 , n345 , n361 , n378 ); 
and ( n380 , n6 , n55 ); 
not ( n381 , n6 ); 
not ( n382 , n148 ); 
and ( n383 , n381 , n382 ); 
nor ( n384 , n380 , n383 ); 
not ( n385 , n384 ); 
and ( n386 , n6 , n186 ); 
not ( n387 , n6 ); 
and ( n388 , n387 , n57 ); 
nor ( n389 , n386 , n388 ); 
not ( n390 , n389 ); 
and ( n391 , n385 , n390 ); 
not ( n392 , n385 ); 
and ( n393 , n392 , n389 ); 
or ( n394 , n391 , n393 ); 
and ( n395 , n6 , n185 ); 
not ( n396 , n6 ); 
and ( n397 , n396 , n60 ); 
nor ( n398 , n395 , n397 ); 
not ( n399 , n398 ); 
not ( n400 , n399 ); 
and ( n401 , n6 , n58 ); 
not ( n402 , n6 ); 
not ( n403 , n147 ); 
and ( n404 , n402 , n403 ); 
nor ( n405 , n401 , n404 ); 
not ( n406 , n405 ); 
not ( n407 , n406 ); 
or ( n408 , n400 , n407 ); 
nand ( n409 , n398 , n405 ); 
nand ( n410 , n408 , n409 ); 
and ( n411 , n394 , n410 ); 
and ( n412 , n6 , n187 ); 
not ( n413 , n6 ); 
and ( n414 , n413 , n54 ); 
nor ( n415 , n412 , n414 ); 
not ( n416 , n415 ); 
not ( n417 , n416 ); 
and ( n418 , n6 , n52 ); 
not ( n419 , n6 ); 
not ( n420 , n149 ); 
and ( n421 , n419 , n420 ); 
nor ( n422 , n418 , n421 ); 
not ( n423 , n422 ); 
not ( n424 , n423 ); 
or ( n425 , n417 , n424 ); 
nand ( n426 , n415 , n422 ); 
nand ( n427 , n425 , n426 ); 
and ( n428 , n6 , n183 ); 
not ( n429 , n6 ); 
and ( n430 , n429 , n66 ); 
nor ( n431 , n428 , n430 ); 
not ( n432 , n64 ); 
and ( n433 , n6 , n432 ); 
not ( n434 , n6 ); 
and ( n435 , n434 , n145 ); 
nor ( n436 , n433 , n435 ); 
nor ( n437 , n431 , n436 ); 
not ( n438 , n437 ); 
nand ( n439 , n431 , n436 ); 
and ( n440 , n6 , n184 ); 
not ( n441 , n6 ); 
and ( n442 , n441 , n63 ); 
nor ( n443 , n440 , n442 ); 
not ( n444 , n443 ); 
not ( n445 , n61 ); 
and ( n446 , n6 , n445 ); 
not ( n447 , n6 ); 
and ( n448 , n447 , n146 ); 
nor ( n449 , n446 , n448 ); 
not ( n450 , n449 ); 
not ( n451 , n450 ); 
or ( n452 , n444 , n451 ); 
not ( n453 , n443 ); 
nand ( n454 , n453 , n449 ); 
nand ( n455 , n452 , n454 ); 
and ( n456 , n427 , n438 , n439 , n455 ); 
and ( n457 , n379 , n411 , n456 ); 
and ( n458 , n6 , n176 ); 
not ( n459 , n6 ); 
and ( n460 , n459 , n29 ); 
nor ( n461 , n458 , n460 ); 
not ( n462 , n461 ); 
and ( n463 , n6 , n28 ); 
not ( n464 , n6 ); 
not ( n465 , n137 ); 
and ( n466 , n464 , n465 ); 
nor ( n467 , n463 , n466 ); 
not ( n468 , n467 ); 
or ( n469 , n462 , n468 ); 
not ( n470 , n461 ); 
not ( n471 , n467 ); 
nand ( n472 , n470 , n471 ); 
nand ( n473 , n469 , n472 ); 
nand ( n474 , n8 , n9 ); 
not ( n475 , n177 ); 
nand ( n476 , n6 , n475 ); 
nand ( n477 , n474 , n476 ); 
not ( n478 , n477 ); 
not ( n479 , n26 ); 
and ( n480 , n6 , n479 ); 
not ( n481 , n6 ); 
and ( n482 , n481 , n138 ); 
nor ( n483 , n480 , n482 ); 
not ( n484 , n483 ); 
not ( n485 , n484 ); 
or ( n486 , n478 , n485 ); 
or ( n487 , n484 , n477 ); 
nand ( n488 , n486 , n487 ); 
and ( n489 , n473 , n488 ); 
not ( n490 , n6 ); 
not ( n491 , n173 ); 
or ( n492 , n490 , n491 ); 
not ( n493 , n6 ); 
nand ( n494 , n493 , n38 ); 
nand ( n495 , n492 , n494 ); 
and ( n496 , n6 , n37 ); 
not ( n497 , n6 ); 
not ( n498 , n134 ); 
and ( n499 , n497 , n498 ); 
nor ( n500 , n496 , n499 ); 
xor ( n501 , n495 , n500 ); 
and ( n502 , n6 , n174 ); 
not ( n503 , n6 ); 
and ( n504 , n503 , n35 ); 
nor ( n505 , n502 , n504 ); 
not ( n506 , n505 ); 
not ( n507 , n34 ); 
and ( n508 , n6 , n507 ); 
not ( n509 , n6 ); 
and ( n510 , n509 , n135 ); 
nor ( n511 , n508 , n510 ); 
not ( n512 , n511 ); 
nand ( n513 , n506 , n512 ); 
nand ( n514 , n505 , n511 ); 
and ( n515 , n6 , n31 ); 
not ( n516 , n6 ); 
not ( n517 , n136 ); 
and ( n518 , n516 , n517 ); 
nor ( n519 , n515 , n518 ); 
not ( n520 , n6 ); 
not ( n521 , n175 ); 
or ( n522 , n520 , n521 ); 
not ( n523 , n6 ); 
nand ( n524 , n523 , n32 ); 
nand ( n525 , n522 , n524 ); 
xor ( n526 , n519 , n525 ); 
nand ( n527 , n513 , n514 , n526 ); 
not ( n528 , n527 ); 
not ( n529 , n168 ); 
nand ( n530 , n6 , n529 ); 
nand ( n531 , n242 , n530 ); 
and ( n532 , n6 , n25 ); 
not ( n533 , n6 ); 
not ( n534 , n128 ); 
and ( n535 , n533 , n534 ); 
nor ( n536 , n532 , n535 ); 
not ( n537 , n536 ); 
and ( n538 , n531 , n537 ); 
not ( n539 , n531 ); 
and ( n540 , n539 , n536 ); 
nor ( n541 , n538 , n540 ); 
nand ( n542 , n8 , n9 ); 
not ( n543 , n169 ); 
nand ( n544 , n6 , n543 ); 
nand ( n545 , n542 , n544 ); 
not ( n546 , n22 ); 
and ( n547 , n6 , n546 ); 
not ( n548 , n6 ); 
and ( n549 , n548 , n129 ); 
nor ( n550 , n547 , n549 ); 
and ( n551 , n545 , n550 ); 
not ( n552 , n545 ); 
not ( n553 , n550 ); 
and ( n554 , n552 , n553 ); 
nor ( n555 , n551 , n554 ); 
nand ( n556 , n541 , n555 ); 
not ( n557 , n171 ); 
nand ( n558 , n6 , n557 ); 
nand ( n559 , n474 , n558 ); 
not ( n560 , n559 ); 
not ( n561 , n560 ); 
and ( n562 , n6 , n18 ); 
not ( n563 , n6 ); 
not ( n564 , n131 ); 
and ( n565 , n563 , n564 ); 
nor ( n566 , n562 , n565 ); 
not ( n567 , n566 ); 
not ( n568 , n567 ); 
or ( n569 , n561 , n568 ); 
nand ( n570 , n559 , n566 ); 
nand ( n571 , n569 , n570 ); 
not ( n572 , n170 ); 
nand ( n573 , n6 , n572 ); 
nand ( n574 , n542 , n573 ); 
not ( n575 , n574 ); 
and ( n576 , n6 , n20 ); 
not ( n577 , n6 ); 
not ( n578 , n130 ); 
and ( n579 , n577 , n578 ); 
nor ( n580 , n576 , n579 ); 
not ( n581 , n580 ); 
or ( n582 , n575 , n581 ); 
or ( n583 , n574 , n580 ); 
nand ( n584 , n582 , n583 ); 
nand ( n585 , n571 , n584 ); 
nor ( n586 , n556 , n585 ); 
and ( n587 , n489 , n501 , n528 , n586 ); 
and ( n588 , n457 , n587 ); 
and ( n589 , n6 , n191 ); 
not ( n590 , n6 ); 
and ( n591 , n590 , n69 ); 
nor ( n592 , n589 , n591 ); 
not ( n593 , n592 ); 
not ( n594 , n67 ); 
and ( n595 , n6 , n594 ); 
not ( n596 , n6 ); 
and ( n597 , n596 , n153 ); 
nor ( n598 , n595 , n597 ); 
not ( n599 , n598 ); 
not ( n600 , n599 ); 
or ( n601 , n593 , n600 ); 
not ( n602 , n592 ); 
nand ( n603 , n602 , n598 ); 
nand ( n604 , n601 , n603 ); 
and ( n605 , n6 , n190 ); 
not ( n606 , n6 ); 
and ( n607 , n606 , n72 ); 
nor ( n608 , n605 , n607 ); 
and ( n609 , n6 , n70 ); 
not ( n610 , n6 ); 
not ( n611 , n152 ); 
and ( n612 , n610 , n611 ); 
nor ( n613 , n609 , n612 ); 
not ( n614 , n613 ); 
xor ( n615 , n608 , n614 ); 
and ( n616 , n6 , n189 ); 
not ( n617 , n6 ); 
and ( n618 , n617 , n75 ); 
nor ( n619 , n616 , n618 ); 
not ( n620 , n619 ); 
and ( n621 , n6 , n73 ); 
not ( n622 , n6 ); 
not ( n623 , n151 ); 
and ( n624 , n622 , n623 ); 
nor ( n625 , n621 , n624 ); 
and ( n626 , n620 , n625 ); 
not ( n627 , n620 ); 
not ( n628 , n625 ); 
and ( n629 , n627 , n628 ); 
nor ( n630 , n626 , n629 ); 
and ( n631 , n6 , n188 ); 
not ( n632 , n6 ); 
and ( n633 , n632 , n77 ); 
nor ( n634 , n631 , n633 ); 
not ( n635 , n634 ); 
and ( n636 , n6 , n78 ); 
not ( n637 , n6 ); 
not ( n638 , n150 ); 
and ( n639 , n637 , n638 ); 
nor ( n640 , n636 , n639 ); 
and ( n641 , n635 , n640 ); 
not ( n642 , n635 ); 
not ( n643 , n640 ); 
and ( n644 , n642 , n643 ); 
nor ( n645 , n641 , n644 ); 
and ( n646 , n604 , n615 , n630 , n645 ); 
not ( n647 , n646 ); 
not ( n648 , n82 ); 
and ( n649 , n6 , n648 ); 
not ( n650 , n6 ); 
and ( n651 , n650 , n159 ); 
nor ( n652 , n649 , n651 ); 
not ( n653 , n652 ); 
and ( n654 , n6 , n196 ); 
not ( n655 , n6 ); 
and ( n656 , n655 , n84 ); 
nor ( n657 , n654 , n656 ); 
not ( n658 , n657 ); 
not ( n659 , n658 ); 
or ( n660 , n653 , n659 ); 
not ( n661 , n652 ); 
nand ( n662 , n657 , n661 ); 
nand ( n663 , n660 , n662 ); 
not ( n664 , n663 ); 
not ( n665 , n88 ); 
and ( n666 , n6 , n665 ); 
not ( n667 , n6 ); 
and ( n668 , n667 , n157 ); 
nor ( n669 , n666 , n668 ); 
nor ( n670 , n664 , n669 ); 
and ( n671 , n6 , n194 ); 
not ( n672 , n6 ); 
and ( n673 , n672 , n90 ); 
nor ( n674 , n671 , n673 ); 
not ( n675 , n674 ); 
and ( n676 , n6 , n197 ); 
not ( n677 , n6 ); 
and ( n678 , n677 , n81 ); 
nor ( n679 , n676 , n678 ); 
not ( n680 , n679 ); 
not ( n681 , n79 ); 
and ( n682 , n6 , n681 ); 
not ( n683 , n6 ); 
and ( n684 , n683 , n160 ); 
nor ( n685 , n682 , n684 ); 
not ( n686 , n685 ); 
xor ( n687 , n680 , n686 ); 
not ( n688 , n687 ); 
and ( n689 , n6 , n195 ); 
not ( n690 , n6 ); 
and ( n691 , n690 , n87 ); 
or ( n692 , n689 , n691 ); 
not ( n693 , n692 ); 
not ( n694 , n85 ); 
and ( n695 , n6 , n694 ); 
not ( n696 , n6 ); 
and ( n697 , n696 , n158 ); 
nor ( n698 , n695 , n697 ); 
not ( n699 , n698 ); 
and ( n700 , n693 , n699 ); 
and ( n701 , n692 , n698 ); 
nor ( n702 , n700 , n701 ); 
nor ( n703 , n688 , n702 ); 
nand ( n704 , n670 , n675 , n703 ); 
and ( n705 , n687 , n661 , n658 ); 
and ( n706 , n680 , n686 ); 
nor ( n707 , n705 , n706 ); 
nand ( n708 , n704 , n707 ); 
not ( n709 , n702 ); 
nand ( n710 , n687 , n709 ); 
not ( n711 , n6 ); 
nand ( n712 , n711 , n156 ); 
not ( n713 , n712 ); 
or ( n714 , n6 , n713 ); 
and ( n715 , n6 , n193 ); 
not ( n716 , n6 ); 
and ( n717 , n716 , n93 ); 
nor ( n718 , n715 , n717 ); 
not ( n719 , n718 ); 
not ( n720 , n6 ); 
nand ( n721 , n719 , n720 ); 
not ( n722 , n721 ); 
nand ( n723 , n714 , n722 ); 
not ( n724 , n723 ); 
and ( n725 , n674 , n669 ); 
not ( n726 , n674 ); 
not ( n727 , n669 ); 
and ( n728 , n726 , n727 ); 
nor ( n729 , n725 , n728 ); 
nand ( n730 , n724 , n663 , n729 ); 
or ( n731 , n710 , n730 ); 
not ( n732 , n692 ); 
nor ( n733 , n732 , n698 ); 
nand ( n734 , n733 , n687 , n663 ); 
nand ( n735 , n731 , n734 ); 
nor ( n736 , n708 , n735 ); 
not ( n737 , n736 ); 
not ( n738 , n737 ); 
or ( n739 , n647 , n738 ); 
nand ( n740 , n640 , n615 ); 
nand ( n741 , n635 , n604 , n630 ); 
or ( n742 , n740 , n741 ); 
or ( n743 , n592 , n598 ); 
nand ( n744 , n742 , n743 ); 
not ( n745 , n604 ); 
or ( n746 , n745 , n614 , n608 ); 
not ( n747 , n628 ); 
nand ( n748 , n620 , n747 , n604 , n615 ); 
nand ( n749 , n746 , n748 ); 
nor ( n750 , n744 , n749 ); 
nand ( n751 , n739 , n750 ); 
nand ( n752 , n588 , n751 ); 
not ( n753 , n714 ); 
nand ( n754 , n753 , n721 ); 
nand ( n755 , n723 , n754 , n729 ); 
nor ( n756 , n755 , n702 ); 
nand ( n757 , n756 , n198 , n687 , n663 ); 
not ( n758 , n757 ); 
and ( n759 , n457 , n587 , n758 , n646 ); 
not ( n760 , n759 ); 
not ( n761 , n586 ); 
not ( n762 , n761 ); 
not ( n763 , n477 ); 
not ( n764 , n763 ); 
not ( n765 , n764 ); 
not ( n766 , n765 ); 
not ( n767 , n484 ); 
or ( n768 , n766 , n767 ); 
buf ( n769 , n467 ); 
not ( n770 , n769 ); 
not ( n771 , n770 ); 
nand ( n772 , n488 , n771 , n470 ); 
nand ( n773 , n768 , n772 ); 
and ( n774 , n519 , n525 ); 
and ( n775 , n473 , n774 , n488 ); 
nor ( n776 , n773 , n775 ); 
not ( n777 , n513 ); 
nand ( n778 , n777 , n473 , n488 , n526 ); 
not ( n779 , n527 ); 
and ( n780 , n495 , n488 ); 
nand ( n781 , n779 , n780 , n500 , n473 ); 
nand ( n782 , n776 , n778 , n781 ); 
nand ( n783 , n762 , n782 ); 
not ( n784 , n574 ); 
nand ( n785 , n580 , n784 , n571 ); 
not ( n786 , n567 ); 
nand ( n787 , n786 , n560 ); 
nand ( n788 , n783 , n785 , n787 ); 
nand ( n789 , n536 , n571 , n584 ); 
buf ( n790 , n531 ); 
not ( n791 , n555 ); 
or ( n792 , n789 , n790 , n791 ); 
nand ( n793 , n571 , n584 ); 
or ( n794 , n793 , n545 , n550 ); 
nand ( n795 , n792 , n794 ); 
nor ( n796 , n788 , n795 ); 
not ( n797 , n379 ); 
buf ( n798 , n384 ); 
nand ( n799 , n798 , n427 ); 
not ( n800 , n389 ); 
not ( n801 , n800 ); 
or ( n802 , n799 , n801 ); 
not ( n803 , n416 ); 
not ( n804 , n803 ); 
not ( n805 , n804 ); 
not ( n806 , n423 ); 
not ( n807 , n806 ); 
or ( n808 , n805 , n807 ); 
nand ( n809 , n802 , n808 ); 
not ( n810 , n809 ); 
and ( n811 , n410 , n455 ); 
nand ( n812 , n811 , n427 , n437 , n394 ); 
buf ( n813 , n449 ); 
not ( n814 , n813 ); 
and ( n815 , n814 , n394 ); 
buf ( n816 , n443 ); 
not ( n817 , n816 ); 
buf ( n818 , n817 ); 
not ( n819 , n427 ); 
not ( n820 , n410 ); 
nor ( n821 , n819 , n820 ); 
nand ( n822 , n815 , n818 , n821 ); 
nand ( n823 , n399 , n405 , n427 , n394 ); 
nand ( n824 , n810 , n812 , n822 , n823 ); 
not ( n825 , n824 ); 
or ( n826 , n797 , n825 ); 
not ( n827 , n320 ); 
not ( n828 , n327 ); 
and ( n829 , n827 , n828 ); 
nor ( n830 , n367 , n344 ); 
and ( n831 , n830 , n373 , n329 , n361 ); 
nor ( n832 , n829 , n831 ); 
not ( n833 , n340 ); 
nand ( n834 , n833 , n335 , n329 ); 
nand ( n835 , n358 , n355 , n329 , n345 ); 
and ( n836 , n832 , n834 , n835 ); 
nand ( n837 , n826 , n836 ); 
nand ( n838 , n837 , n587 ); 
nand ( n839 , n752 , n760 , n796 , n838 ); 
not ( n840 , n839 ); 
or ( n841 , n315 , n840 ); 
not ( n842 , n236 ); 
not ( n843 , n246 ); 
not ( n844 , n285 ); 
or ( n845 , n842 , n843 , n844 ); 
or ( n846 , n273 , n281 ); 
nand ( n847 , n845 , n846 ); 
not ( n848 , n312 ); 
nand ( n849 , n267 , n848 ); 
not ( n850 , n293 ); 
nand ( n851 , n285 , n850 , n248 ); 
nor ( n852 , n849 , n851 ); 
nor ( n853 , n847 , n852 ); 
nand ( n854 , n256 , n262 , n285 , n248 ); 
not ( n855 , n267 ); 
nor ( n856 , n301 , n855 ); 
nand ( n857 , n856 , n308 , n285 , n248 ); 
nand ( n858 , n853 , n854 , n857 ); 
not ( n859 , n858 ); 
nand ( n860 , n841 , n859 ); 
not ( n861 , n225 ); 
xnor ( n862 , n3 , n219 ); 
nor ( n863 , n861 , n862 ); 
nand ( n864 , n860 , n863 ); 
nand ( n865 , n229 , n864 ); 
nand ( n866 , n863 , n858 ); 
and ( n867 , n863 , n314 ); 
nand ( n868 , n867 , n759 ); 
nand ( n869 , n867 , n588 , n751 ); 
and ( n870 , n866 , n868 , n869 ); 
nand ( n871 , n796 , n838 ); 
nand ( n872 , n867 , n871 ); 
nand ( n873 , n870 , n229 , n872 ); 
not ( n874 , n10 ); 
not ( n875 , n874 ); 
not ( n876 , n6 ); 
not ( n877 , n11 ); 
not ( n878 , n877 ); 
or ( n879 , n876 , n878 ); 
nand ( n880 , n879 , n242 ); 
not ( n881 , n880 ); 
not ( n882 , n881 ); 
not ( n883 , n882 ); 
or ( n884 , n875 , n883 ); 
not ( n885 , n881 ); 
or ( n886 , n885 , n874 ); 
nand ( n887 , n884 , n886 ); 
not ( n888 , n887 ); 
nand ( n889 , n1 , n4 ); 
or ( n890 , n3 , n889 ); 
nand ( n891 , n3 , n889 ); 
nand ( n892 , n1 , n2 ); 
and ( n893 , n892 , n3 ); 
not ( n894 , n892 ); 
and ( n895 , n894 , n223 ); 
nor ( n896 , n893 , n895 ); 
nand ( n897 , n890 , n891 , n896 ); 
nor ( n898 , n888 , n897 ); 
not ( n899 , n5 ); 
not ( n900 , n7 ); 
nand ( n901 , n6 , n900 ); 
nand ( n902 , n242 , n901 ); 
not ( n903 , n902 ); 
not ( n904 , n903 ); 
and ( n905 , n899 , n904 ); 
and ( n906 , n5 , n903 ); 
nor ( n907 , n905 , n906 ); 
not ( n908 , n907 ); 
not ( n909 , n908 ); 
not ( n910 , n909 ); 
not ( n911 , n303 ); 
not ( n912 , n15 ); 
nand ( n913 , n912 , n6 ); 
nand ( n914 , n913 , n254 ); 
not ( n915 , n914 ); 
or ( n916 , n911 , n915 ); 
or ( n917 , n303 , n914 ); 
nand ( n918 , n916 , n917 ); 
not ( n919 , n17 ); 
nand ( n920 , n6 , n919 ); 
nand ( n921 , n254 , n920 ); 
and ( n922 , n16 , n921 ); 
nor ( n923 , n16 , n921 ); 
not ( n924 , n13 ); 
nand ( n925 , n6 , n924 ); 
nand ( n926 , n254 , n925 ); 
not ( n927 , n12 ); 
and ( n928 , n926 , n927 ); 
not ( n929 , n926 ); 
and ( n930 , n929 , n12 ); 
nor ( n931 , n928 , n930 ); 
nor ( n932 , n922 , n923 , n931 ); 
and ( n933 , n898 , n910 , n918 , n932 ); 
not ( n934 , n52 ); 
and ( n935 , n6 , n53 ); 
not ( n936 , n6 ); 
and ( n937 , n936 , n54 ); 
nor ( n938 , n935 , n937 ); 
not ( n939 , n938 ); 
not ( n940 , n939 ); 
or ( n941 , n934 , n940 ); 
not ( n942 , n52 ); 
nand ( n943 , n942 , n938 ); 
nand ( n944 , n941 , n943 ); 
not ( n945 , n58 ); 
and ( n946 , n6 , n59 ); 
not ( n947 , n6 ); 
and ( n948 , n947 , n60 ); 
nor ( n949 , n946 , n948 ); 
not ( n950 , n949 ); 
not ( n951 , n950 ); 
and ( n952 , n945 , n951 ); 
and ( n953 , n58 , n950 ); 
nor ( n954 , n952 , n953 ); 
not ( n955 , n954 ); 
and ( n956 , n944 , n955 ); 
and ( n957 , n6 , n65 ); 
not ( n958 , n6 ); 
and ( n959 , n958 , n66 ); 
or ( n960 , n957 , n959 ); 
xor ( n961 , n432 , n960 ); 
and ( n962 , n6 , n41 ); 
not ( n963 , n6 ); 
and ( n964 , n963 , n42 ); 
nor ( n965 , n962 , n964 ); 
and ( n966 , n965 , n40 ); 
not ( n967 , n965 ); 
not ( n968 , n40 ); 
and ( n969 , n967 , n968 ); 
or ( n970 , n966 , n969 ); 
and ( n971 , n6 , n47 ); 
not ( n972 , n6 ); 
and ( n973 , n972 , n48 ); 
nor ( n974 , n971 , n973 ); 
xnor ( n975 , n974 , n46 ); 
nor ( n976 , n970 , n975 ); 
and ( n977 , n6 , n44 ); 
not ( n978 , n6 ); 
and ( n979 , n978 , n45 ); 
or ( n980 , n977 , n979 ); 
and ( n981 , n980 , n330 ); 
not ( n982 , n980 ); 
and ( n983 , n982 , n43 ); 
nor ( n984 , n981 , n983 ); 
not ( n985 , n51 ); 
not ( n986 , n6 ); 
not ( n987 , n49 ); 
or ( n988 , n986 , n987 ); 
nand ( n989 , n988 , n372 ); 
not ( n990 , n989 ); 
or ( n991 , n985 , n990 ); 
or ( n992 , n51 , n989 ); 
nand ( n993 , n991 , n992 ); 
and ( n994 , n984 , n993 ); 
and ( n995 , n956 , n961 , n976 , n994 ); 
not ( n996 , n55 ); 
and ( n997 , n6 , n56 ); 
not ( n998 , n6 ); 
and ( n999 , n998 , n57 ); 
nor ( n1000 , n997 , n999 ); 
not ( n1001 , n1000 ); 
not ( n1002 , n1001 ); 
and ( n1003 , n996 , n1002 ); 
and ( n1004 , n55 , n1001 ); 
nor ( n1005 , n1003 , n1004 ); 
not ( n1006 , n1005 ); 
and ( n1007 , n6 , n62 ); 
not ( n1008 , n6 ); 
and ( n1009 , n1008 , n63 ); 
nor ( n1010 , n1007 , n1009 ); 
and ( n1011 , n1010 , n445 ); 
not ( n1012 , n1010 ); 
and ( n1013 , n1012 , n61 ); 
nor ( n1014 , n1011 , n1013 ); 
not ( n1015 , n1014 ); 
and ( n1016 , n995 , n1006 , n1015 ); 
and ( n1017 , n933 , n1016 ); 
and ( n1018 , n6 , n68 ); 
not ( n1019 , n6 ); 
and ( n1020 , n1019 , n69 ); 
nor ( n1021 , n1018 , n1020 ); 
and ( n1022 , n1021 , n67 ); 
not ( n1023 , n1021 ); 
and ( n1024 , n1023 , n594 ); 
nor ( n1025 , n1022 , n1024 ); 
not ( n1026 , n1025 ); 
and ( n1027 , n6 , n71 ); 
not ( n1028 , n6 ); 
and ( n1029 , n1028 , n72 ); 
nor ( n1030 , n1027 , n1029 ); 
not ( n1031 , n1030 ); 
and ( n1032 , n70 , n1031 ); 
not ( n1033 , n70 ); 
and ( n1034 , n1033 , n1030 ); 
nor ( n1035 , n1032 , n1034 ); 
and ( n1036 , n6 , n76 ); 
not ( n1037 , n6 ); 
and ( n1038 , n1037 , n77 ); 
nor ( n1039 , n1036 , n1038 ); 
not ( n1040 , n1039 ); 
and ( n1041 , n78 , n1040 ); 
nor ( n1042 , n78 , n1040 ); 
nor ( n1043 , n1041 , n1042 ); 
and ( n1044 , n6 , n74 ); 
not ( n1045 , n6 ); 
and ( n1046 , n1045 , n75 ); 
nor ( n1047 , n1044 , n1046 ); 
xnor ( n1048 , n1047 , n73 ); 
nor ( n1049 , n1026 , n1035 , n1043 , n1048 ); 
and ( n1050 , n6 , n92 ); 
not ( n1051 , n6 ); 
and ( n1052 , n1051 , n93 ); 
nor ( n1053 , n1050 , n1052 ); 
not ( n1054 , n1053 ); 
nand ( n1055 , n1054 , n720 ); 
not ( n1056 , n6 ); 
nand ( n1057 , n1056 , n91 ); 
not ( n1058 , n1057 ); 
and ( n1059 , n1055 , n1058 ); 
not ( n1060 , n1055 ); 
and ( n1061 , n1060 , n1057 ); 
nor ( n1062 , n1059 , n1061 ); 
and ( n1063 , n6 , n80 ); 
not ( n1064 , n6 ); 
and ( n1065 , n1064 , n81 ); 
nor ( n1066 , n1063 , n1065 ); 
not ( n1067 , n1066 ); 
xor ( n1068 , n681 , n1067 ); 
and ( n1069 , n6 , n86 ); 
not ( n1070 , n6 ); 
and ( n1071 , n1070 , n87 ); 
nor ( n1072 , n1069 , n1071 ); 
and ( n1073 , n694 , n1072 ); 
not ( n1074 , n694 ); 
not ( n1075 , n1072 ); 
and ( n1076 , n1074 , n1075 ); 
nor ( n1077 , n1073 , n1076 ); 
not ( n1078 , n1077 ); 
nand ( n1079 , n94 , n1062 , n1068 , n1078 ); 
and ( n1080 , n6 , n83 ); 
not ( n1081 , n6 ); 
and ( n1082 , n1081 , n84 ); 
nor ( n1083 , n1080 , n1082 ); 
and ( n1084 , n1083 , n82 ); 
not ( n1085 , n1083 ); 
not ( n1086 , n82 ); 
and ( n1087 , n1085 , n1086 ); 
or ( n1088 , n1084 , n1087 ); 
and ( n1089 , n6 , n89 ); 
not ( n1090 , n6 ); 
and ( n1091 , n1090 , n90 ); 
nor ( n1092 , n1089 , n1091 ); 
and ( n1093 , n1092 , n665 ); 
not ( n1094 , n1092 ); 
and ( n1095 , n1094 , n88 ); 
nor ( n1096 , n1093 , n1095 ); 
nor ( n1097 , n1079 , n1088 , n1096 ); 
and ( n1098 , n6 , n30 ); 
not ( n1099 , n6 ); 
and ( n1100 , n1099 , n29 ); 
nor ( n1101 , n1098 , n1100 ); 
and ( n1102 , n28 , n1101 ); 
not ( n1103 , n1102 ); 
not ( n1104 , n28 ); 
not ( n1105 , n1101 ); 
nand ( n1106 , n1104 , n1105 ); 
nand ( n1107 , n1103 , n1106 ); 
not ( n1108 , n1107 ); 
not ( n1109 , n1108 ); 
not ( n1110 , n1109 ); 
and ( n1111 , n6 , n36 ); 
not ( n1112 , n6 ); 
and ( n1113 , n1112 , n35 ); 
nor ( n1114 , n1111 , n1113 ); 
and ( n1115 , n1114 , n34 ); 
not ( n1116 , n1114 ); 
and ( n1117 , n1116 , n507 ); 
nor ( n1118 , n1115 , n1117 ); 
not ( n1119 , n1118 ); 
nor ( n1120 , n1110 , n1119 ); 
and ( n1121 , n6 , n39 ); 
not ( n1122 , n6 ); 
and ( n1123 , n1122 , n38 ); 
nor ( n1124 , n1121 , n1123 ); 
not ( n1125 , n1124 ); 
and ( n1126 , n37 , n1125 ); 
nor ( n1127 , n37 , n1125 ); 
nor ( n1128 , n1126 , n1127 ); 
not ( n1129 , n6 ); 
not ( n1130 , n21 ); 
not ( n1131 , n1130 ); 
or ( n1132 , n1129 , n1131 ); 
nand ( n1133 , n1132 , n254 ); 
not ( n1134 , n1133 ); 
and ( n1135 , n20 , n1134 ); 
not ( n1136 , n20 ); 
and ( n1137 , n1136 , n1133 ); 
or ( n1138 , n1135 , n1137 ); 
not ( n1139 , n24 ); 
nand ( n1140 , n6 , n1139 ); 
nand ( n1141 , n254 , n1140 ); 
and ( n1142 , n1141 , n25 ); 
not ( n1143 , n1141 ); 
not ( n1144 , n25 ); 
and ( n1145 , n1143 , n1144 ); 
nor ( n1146 , n1142 , n1145 ); 
not ( n1147 , n23 ); 
nand ( n1148 , n6 , n1147 ); 
nand ( n1149 , n254 , n1148 ); 
and ( n1150 , n1149 , n22 ); 
not ( n1151 , n1149 ); 
and ( n1152 , n1151 , n546 ); 
nor ( n1153 , n1150 , n1152 ); 
not ( n1154 , n18 ); 
buf ( n1155 , n6 ); 
buf ( n1156 , n6 ); 
nand ( n1157 , n6 , n1156 , n19 ); 
nand ( n1158 , n1155 , n242 , n1157 ); 
not ( n1159 , n1158 ); 
not ( n1160 , n1159 ); 
or ( n1161 , n1154 , n1160 ); 
not ( n1162 , n1158 ); 
or ( n1163 , n18 , n1162 ); 
nand ( n1164 , n1161 , n1163 ); 
nand ( n1165 , n1138 , n1146 , n1153 , n1164 ); 
nor ( n1166 , n1128 , n1165 ); 
not ( n1167 , n31 ); 
not ( n1168 , n6 ); 
not ( n1169 , n33 ); 
or ( n1170 , n1168 , n1169 ); 
nand ( n1171 , n1170 , n524 ); 
xor ( n1172 , n1167 , n1171 ); 
not ( n1173 , n6 ); 
nand ( n1174 , n6 , n27 ); 
nor ( n1175 , n1173 , n1174 ); 
not ( n1176 , n1175 ); 
not ( n1177 , n6 ); 
nand ( n1178 , n1177 , n1174 ); 
nand ( n1179 , n1176 , n242 , n1178 ); 
not ( n1180 , n1179 ); 
and ( n1181 , n1180 , n26 ); 
not ( n1182 , n1180 ); 
not ( n1183 , n26 ); 
and ( n1184 , n1182 , n1183 ); 
nor ( n1185 , n1181 , n1184 ); 
not ( n1186 , n1185 ); 
and ( n1187 , n1120 , n1166 , n1172 , n1186 ); 
nand ( n1188 , n1017 , n1049 , n1097 , n1187 ); 
nor ( n1189 , n78 , n1035 , n1048 ); 
and ( n1190 , n1189 , n1040 , n1025 ); 
not ( n1191 , n1025 ); 
nor ( n1192 , n1191 , n73 , n1047 , n1035 ); 
nor ( n1193 , n1190 , n1192 ); 
not ( n1194 , n1021 ); 
nand ( n1195 , n1194 , n594 ); 
not ( n1196 , n70 ); 
nand ( n1197 , n1196 , n1031 , n1025 ); 
not ( n1198 , n1088 ); 
nor ( n1199 , n85 , n1072 ); 
nand ( n1200 , n1198 , n1199 , n1068 ); 
not ( n1201 , n88 ); 
not ( n1202 , n1092 ); 
not ( n1203 , n1202 ); 
nor ( n1204 , n1203 , n1088 ); 
nand ( n1205 , n1201 , n1204 , n1068 , n1078 ); 
not ( n1206 , n1083 ); 
and ( n1207 , n1086 , n1206 , n1068 ); 
and ( n1208 , n681 , n1067 ); 
nor ( n1209 , n1207 , n1208 ); 
nor ( n1210 , n1055 , n1088 ); 
nor ( n1211 , n1077 , n1096 ); 
nand ( n1212 , n1210 , n1211 , n1057 , n1068 ); 
nand ( n1213 , n1200 , n1205 , n1209 , n1212 ); 
nand ( n1214 , n1049 , n1213 ); 
nand ( n1215 , n1193 , n1195 , n1197 , n1214 ); 
nand ( n1216 , n933 , n1016 , n1187 , n1215 ); 
nand ( n1217 , n3 , n892 ); 
not ( n1218 , n896 ); 
nor ( n1219 , n1218 , n891 ); 
and ( n1220 , n1217 , n1219 ); 
nor ( n1221 , n1217 , n1219 ); 
or ( n1222 , n10 , n885 , n907 ); 
or ( n1223 , n5 , n902 ); 
nand ( n1224 , n1222 , n1223 ); 
not ( n1225 , n887 ); 
nor ( n1226 , n1225 , n12 , n926 , n907 ); 
nor ( n1227 , n1224 , n1226 ); 
and ( n1228 , n908 , n923 , n918 ); 
not ( n1229 , n931 ); 
and ( n1230 , n1228 , n887 , n1229 ); 
nor ( n1231 , n914 , n909 ); 
nand ( n1232 , n887 , n1229 ); 
nor ( n1233 , n14 , n1232 ); 
and ( n1234 , n1231 , n1233 ); 
nor ( n1235 , n1230 , n1234 ); 
and ( n1236 , n1227 , n1235 ); 
nor ( n1237 , n1236 , n897 ); 
nor ( n1238 , n1220 , n1221 , n1237 ); 
not ( n1239 , n1187 ); 
nor ( n1240 , n51 , n970 , n975 ); 
and ( n1241 , n1240 , n989 , n984 ); 
not ( n1242 , n984 ); 
nor ( n1243 , n1242 , n46 , n974 , n970 ); 
nor ( n1244 , n1241 , n1243 ); 
not ( n1245 , n965 ); 
nand ( n1246 , n1245 , n968 ); 
not ( n1247 , n43 ); 
not ( n1248 , n970 ); 
nand ( n1249 , n1247 , n980 , n1248 ); 
nand ( n1250 , n976 , n994 ); 
not ( n1251 , n1250 ); 
not ( n1252 , n942 ); 
not ( n1253 , n939 ); 
or ( n1254 , n1252 , n1253 ); 
not ( n1255 , n55 ); 
nand ( n1256 , n1255 , n1001 , n944 ); 
nand ( n1257 , n1254 , n1256 ); 
not ( n1258 , n1257 ); 
not ( n1259 , n58 ); 
nand ( n1260 , n1259 , n944 , n1006 , n950 ); 
not ( n1261 , n1010 ); 
not ( n1262 , n1261 ); 
not ( n1263 , n944 ); 
nor ( n1264 , n1262 , n1263 ); 
nand ( n1265 , n1264 , n445 , n1006 , n955 ); 
and ( n1266 , n432 , n960 ); 
nor ( n1267 , n1263 , n954 ); 
nor ( n1268 , n1005 , n1014 ); 
nand ( n1269 , n1266 , n1267 , n1268 ); 
nand ( n1270 , n1258 , n1260 , n1265 , n1269 ); 
nand ( n1271 , n1251 , n1270 ); 
nand ( n1272 , n1244 , n1246 , n1249 , n1271 ); 
not ( n1273 , n1272 ); 
or ( n1274 , n1239 , n1273 ); 
not ( n1275 , n1153 ); 
not ( n1276 , n1164 ); 
nor ( n1277 , n25 , n1275 , n1276 ); 
not ( n1278 , n1141 ); 
and ( n1279 , n1277 , n1278 , n1138 ); 
not ( n1280 , n1138 ); 
buf ( n1281 , n1149 ); 
nor ( n1282 , n1280 , n22 , n1281 , n1276 ); 
nor ( n1283 , n1279 , n1282 ); 
not ( n1284 , n18 ); 
nand ( n1285 , n1284 , n1162 ); 
not ( n1286 , n20 ); 
not ( n1287 , n1276 ); 
nand ( n1288 , n1286 , n1134 , n1287 ); 
not ( n1289 , n1165 ); 
and ( n1290 , n1167 , n1171 ); 
nor ( n1291 , n1108 , n1185 ); 
and ( n1292 , n1290 , n1291 ); 
or ( n1293 , n1106 , n1185 ); 
buf ( n1294 , n1179 ); 
not ( n1295 , n1294 ); 
not ( n1296 , n1295 ); 
or ( n1297 , n26 , n1296 ); 
nand ( n1298 , n1293 , n1297 ); 
nor ( n1299 , n1292 , n1298 ); 
not ( n1300 , n1114 ); 
and ( n1301 , n1300 , n1172 ); 
nand ( n1302 , n1301 , n507 , n1109 , n1186 ); 
nor ( n1303 , n37 , n1124 ); 
and ( n1304 , n1172 , n1118 ); 
not ( n1305 , n1185 ); 
nand ( n1306 , n1303 , n1304 , n1109 , n1305 ); 
nand ( n1307 , n1299 , n1302 , n1306 ); 
nand ( n1308 , n1289 , n1307 ); 
and ( n1309 , n1283 , n1285 , n1288 , n1308 ); 
nand ( n1310 , n1274 , n1309 ); 
nand ( n1311 , n933 , n1310 ); 
nand ( n1312 , n1188 , n1216 , n1238 , n1311 ); 
not ( n1313 , n824 ); 
not ( n1314 , n1313 ); 
not ( n1315 , n750 ); 
not ( n1316 , n757 ); 
not ( n1317 , n736 ); 
or ( n1318 , n1316 , n1317 ); 
nand ( n1319 , n1318 , n646 ); 
not ( n1320 , n1319 ); 
or ( n1321 , n1315 , n1320 ); 
and ( n1322 , n411 , n456 ); 
nand ( n1323 , n1321 , n1322 ); 
not ( n1324 , n1323 ); 
or ( n1325 , n1314 , n1324 ); 
nand ( n1326 , n1325 , n379 ); 
nand ( n1327 , n836 , n1326 ); 
not ( n1328 , n620 ); 
not ( n1329 , n634 ); 
or ( n1330 , n1328 , n1329 ); 
nand ( n1331 , n635 , n619 ); 
nand ( n1332 , n1330 , n1331 ); 
and ( n1333 , n608 , n602 ); 
not ( n1334 , n608 ); 
and ( n1335 , n1334 , n592 ); 
or ( n1336 , n1333 , n1335 ); 
xor ( n1337 , n1332 , n1336 ); 
and ( n1338 , n679 , n658 ); 
not ( n1339 , n679 ); 
and ( n1340 , n1339 , n657 ); 
or ( n1341 , n1338 , n1340 ); 
not ( n1342 , n6 ); 
not ( n1343 , n192 ); 
or ( n1344 , n1342 , n1343 ); 
not ( n1345 , n6 ); 
nand ( n1346 , n1345 , n118 ); 
nand ( n1347 , n1344 , n1346 ); 
not ( n1348 , n1347 ); 
not ( n1349 , n718 ); 
or ( n1350 , n1348 , n1349 ); 
or ( n1351 , n718 , n1347 ); 
nand ( n1352 , n1350 , n1351 ); 
not ( n1353 , n1352 ); 
and ( n1354 , n1341 , n1353 ); 
not ( n1355 , n1341 ); 
and ( n1356 , n1355 , n1352 ); 
nor ( n1357 , n1354 , n1356 ); 
not ( n1358 , n675 ); 
not ( n1359 , n732 ); 
or ( n1360 , n1358 , n1359 ); 
nand ( n1361 , n692 , n674 ); 
nand ( n1362 , n1360 , n1361 ); 
not ( n1363 , n1362 ); 
and ( n1364 , n1357 , n1363 ); 
not ( n1365 , n1357 ); 
and ( n1366 , n1365 , n1362 ); 
nor ( n1367 , n1364 , n1366 ); 
not ( n1368 , n1367 ); 
and ( n1369 , n1337 , n1368 ); 
not ( n1370 , n1337 ); 
and ( n1371 , n1370 , n1367 ); 
nor ( n1372 , n1369 , n1371 ); 
not ( n1373 , n833 ); 
not ( n1374 , n320 ); 
or ( n1375 , n1373 , n1374 ); 
nand ( n1376 , n319 , n340 ); 
nand ( n1377 , n1375 , n1376 ); 
not ( n1378 , n358 ); 
not ( n1379 , n374 ); 
or ( n1380 , n1378 , n1379 ); 
nand ( n1381 , n373 , n349 ); 
nand ( n1382 , n1380 , n1381 ); 
xnor ( n1383 , n1377 , n1382 ); 
not ( n1384 , n804 ); 
not ( n1385 , n800 ); 
not ( n1386 , n1385 ); 
or ( n1387 , n1384 , n1386 ); 
nand ( n1388 , n800 , n803 ); 
nand ( n1389 , n1387 , n1388 ); 
and ( n1390 , n6 , n182 ); 
not ( n1391 , n6 ); 
and ( n1392 , n1391 , n116 ); 
or ( n1393 , n1390 , n1392 ); 
not ( n1394 , n1393 ); 
not ( n1395 , n431 ); 
or ( n1396 , n1394 , n1395 ); 
or ( n1397 , n431 , n1393 ); 
nand ( n1398 , n1396 , n1397 ); 
not ( n1399 , n1398 ); 
and ( n1400 , n1389 , n1399 ); 
not ( n1401 , n1389 ); 
and ( n1402 , n1401 , n1398 ); 
nor ( n1403 , n1400 , n1402 ); 
and ( n1404 , n399 , n817 ); 
not ( n1405 , n399 ); 
and ( n1406 , n1405 , n816 ); 
nor ( n1407 , n1404 , n1406 ); 
and ( n1408 , n1403 , n1407 ); 
not ( n1409 , n1403 ); 
not ( n1410 , n1407 ); 
and ( n1411 , n1409 , n1410 ); 
nor ( n1412 , n1408 , n1411 ); 
not ( n1413 , n1412 ); 
and ( n1414 , n1383 , n1413 ); 
not ( n1415 , n1383 ); 
and ( n1416 , n1415 , n1412 ); 
nor ( n1417 , n1414 , n1416 ); 
nor ( n1418 , n1372 , n1417 ); 
not ( n1419 , n301 ); 
not ( n1420 , n256 ); 
or ( n1421 , n1419 , n1420 ); 
not ( n1422 , n301 ); 
nand ( n1423 , n1422 , n255 ); 
nand ( n1424 , n1421 , n1423 ); 
not ( n1425 , n1424 ); 
not ( n1426 , n243 ); 
not ( n1427 , n274 ); 
or ( n1428 , n1426 , n1427 ); 
not ( n1429 , n243 ); 
nand ( n1430 , n1429 , n273 ); 
nand ( n1431 , n1428 , n1430 ); 
not ( n1432 , n163 ); 
nand ( n1433 , n6 , n1432 ); 
nand ( n1434 , n254 , n1433 ); 
not ( n1435 , n254 ); 
not ( n1436 , n1435 ); 
and ( n1437 , n1434 , n1436 ); 
nor ( n1438 , n1437 , 1'b0 ); 
not ( n1439 , n1438 ); 
and ( n1440 , n1431 , n1439 ); 
not ( n1441 , n1431 ); 
and ( n1442 , n1441 , n1438 ); 
nor ( n1443 , n1440 , n1442 ); 
not ( n1444 , n1443 ); 
or ( n1445 , n1425 , n1444 ); 
or ( n1446 , n1424 , n1443 ); 
nand ( n1447 , n1445 , n1446 ); 
xor ( n1448 , n162 , n161 ); 
and ( n1449 , n1448 , n287 , n6 ); 
and ( n1450 , n1447 , n1449 ); 
not ( n1451 , n1447 ); 
not ( n1452 , n1449 ); 
and ( n1453 , n1451 , n1452 ); 
nor ( n1454 , n1450 , n1453 ); 
not ( n1455 , n790 ); 
and ( n1456 , n545 , n1455 ); 
not ( n1457 , n545 ); 
and ( n1458 , n1457 , n790 ); 
nor ( n1459 , n1456 , n1458 ); 
not ( n1460 , n1459 ); 
or ( n1461 , n784 , n559 ); 
or ( n1462 , n560 , n574 ); 
nand ( n1463 , n1461 , n1462 ); 
not ( n1464 , n1463 ); 
and ( n1465 , n1460 , n1464 ); 
and ( n1466 , n1463 , n1459 ); 
nor ( n1467 , n1465 , n1466 ); 
not ( n1468 , n1467 ); 
not ( n1469 , n525 ); 
not ( n1470 , n505 ); 
or ( n1471 , n1469 , n1470 ); 
or ( n1472 , n505 , n525 ); 
nand ( n1473 , n1471 , n1472 ); 
not ( n1474 , n1473 ); 
not ( n1475 , n470 ); 
not ( n1476 , n764 ); 
or ( n1477 , n1475 , n1476 ); 
nand ( n1478 , n461 , n763 ); 
nand ( n1479 , n1477 , n1478 ); 
and ( n1480 , n6 , n172 ); 
not ( n1481 , n6 ); 
and ( n1482 , n1481 , n113 ); 
nor ( n1483 , n1480 , n1482 ); 
not ( n1484 , n1483 ); 
not ( n1485 , n495 ); 
and ( n1486 , n1484 , n1485 ); 
and ( n1487 , n495 , n1483 ); 
nor ( n1488 , n1486 , n1487 ); 
and ( n1489 , n1479 , n1488 ); 
not ( n1490 , n1479 ); 
not ( n1491 , n1488 ); 
and ( n1492 , n1490 , n1491 ); 
nor ( n1493 , n1489 , n1492 ); 
not ( n1494 , n1493 ); 
or ( n1495 , n1474 , n1494 ); 
or ( n1496 , n1473 , n1493 ); 
nand ( n1497 , n1495 , n1496 ); 
not ( n1498 , n1497 ); 
or ( n1499 , n1468 , n1498 ); 
or ( n1500 , n1467 , n1497 ); 
nand ( n1501 , n1499 , n1500 ); 
nand ( n1502 , n1418 , n1454 , n1501 ); 
not ( n1503 , n1502 ); 
xor ( n1504 , n965 , n980 ); 
not ( n1505 , n1504 ); 
xnor ( n1506 , n974 , n989 ); 
not ( n1507 , n1506 ); 
and ( n1508 , n1505 , n1507 ); 
and ( n1509 , n1506 , n1504 ); 
nor ( n1510 , n1508 , n1509 ); 
not ( n1511 , n939 ); 
not ( n1512 , n1000 ); 
or ( n1513 , n1511 , n1512 ); 
nand ( n1514 , n1001 , n938 ); 
nand ( n1515 , n1513 , n1514 ); 
not ( n1516 , n960 ); 
and ( n1517 , n6 , n115 ); 
not ( n1518 , n6 ); 
and ( n1519 , n1518 , n116 ); 
nor ( n1520 , n1517 , n1519 ); 
not ( n1521 , n1520 ); 
or ( n1522 , n1516 , n1521 ); 
or ( n1523 , n1520 , n960 ); 
nand ( n1524 , n1522 , n1523 ); 
not ( n1525 , n1524 ); 
and ( n1526 , n1515 , n1525 ); 
not ( n1527 , n1515 ); 
and ( n1528 , n1527 , n1524 ); 
nor ( n1529 , n1526 , n1528 ); 
not ( n1530 , n950 ); 
not ( n1531 , n1262 ); 
or ( n1532 , n1530 , n1531 ); 
nand ( n1533 , n1261 , n949 ); 
nand ( n1534 , n1532 , n1533 ); 
and ( n1535 , n1529 , n1534 ); 
not ( n1536 , n1529 ); 
not ( n1537 , n1534 ); 
and ( n1538 , n1536 , n1537 ); 
nor ( n1539 , n1535 , n1538 ); 
not ( n1540 , n1539 ); 
and ( n1541 , n1510 , n1540 ); 
not ( n1542 , n1510 ); 
and ( n1543 , n1542 , n1539 ); 
nor ( n1544 , n1541 , n1543 ); 
and ( n1545 , n1021 , n1031 ); 
not ( n1546 , n1021 ); 
and ( n1547 , n1546 , n1030 ); 
nor ( n1548 , n1545 , n1547 ); 
not ( n1549 , n1548 ); 
and ( n1550 , n1047 , n1039 ); 
not ( n1551 , n1047 ); 
and ( n1552 , n1551 , n1040 ); 
nor ( n1553 , n1550 , n1552 ); 
not ( n1554 , n1553 ); 
and ( n1555 , n1549 , n1554 ); 
and ( n1556 , n1553 , n1548 ); 
nor ( n1557 , n1555 , n1556 ); 
not ( n1558 , n1067 ); 
not ( n1559 , n1083 ); 
or ( n1560 , n1558 , n1559 ); 
nand ( n1561 , n1206 , n1066 ); 
nand ( n1562 , n1560 , n1561 ); 
not ( n1563 , n6 ); 
not ( n1564 , n117 ); 
or ( n1565 , n1563 , n1564 ); 
nand ( n1566 , n1565 , n1346 ); 
not ( n1567 , n1566 ); 
not ( n1568 , n1053 ); 
or ( n1569 , n1567 , n1568 ); 
or ( n1570 , n1053 , n1566 ); 
nand ( n1571 , n1569 , n1570 ); 
and ( n1572 , n1562 , n1571 ); 
not ( n1573 , n1562 ); 
not ( n1574 , n1571 ); 
and ( n1575 , n1573 , n1574 ); 
nor ( n1576 , n1572 , n1575 ); 
not ( n1577 , n1075 ); 
not ( n1578 , n1203 ); 
or ( n1579 , n1577 , n1578 ); 
nand ( n1580 , n1202 , n1072 ); 
nand ( n1581 , n1579 , n1580 ); 
and ( n1582 , n1576 , n1581 ); 
not ( n1583 , n1576 ); 
not ( n1584 , n1581 ); 
and ( n1585 , n1583 , n1584 ); 
nor ( n1586 , n1582 , n1585 ); 
and ( n1587 , n1557 , n1586 ); 
not ( n1588 , n1557 ); 
not ( n1589 , n1586 ); 
and ( n1590 , n1588 , n1589 ); 
nor ( n1591 , n1587 , n1590 ); 
nor ( n1592 , n1544 , n1591 ); 
xor ( n1593 , n112 , n111 ); 
and ( n1594 , n1593 , n287 , n6 ); 
not ( n1595 , n1594 ); 
not ( n1596 , n880 ); 
not ( n1597 , n903 ); 
or ( n1598 , n1596 , n1597 ); 
not ( n1599 , n880 ); 
nand ( n1600 , n1599 , n902 ); 
nand ( n1601 , n1598 , n1600 ); 
not ( n1602 , n1435 ); 
not ( n1603 , n921 ); 
and ( n1604 , n1602 , n1603 ); 
not ( n1605 , n1602 ); 
and ( n1606 , n1605 , n921 ); 
nor ( n1607 , n1604 , n1606 ); 
not ( n1608 , n1607 ); 
and ( n1609 , n1601 , n1608 ); 
not ( n1610 , n1601 ); 
and ( n1611 , n1610 , n1607 ); 
nor ( n1612 , n1609 , n1611 ); 
and ( n1613 , n914 , n926 ); 
not ( n1614 , n914 ); 
not ( n1615 , n926 ); 
and ( n1616 , n1614 , n1615 ); 
nor ( n1617 , n1613 , n1616 ); 
not ( n1618 , n1617 ); 
and ( n1619 , n1612 , n1618 ); 
not ( n1620 , n1612 ); 
and ( n1621 , n1620 , n1617 ); 
nor ( n1622 , n1619 , n1621 ); 
not ( n1623 , n1622 ); 
or ( n1624 , n1595 , n1623 ); 
or ( n1625 , n1594 , n1622 ); 
nand ( n1626 , n1624 , n1625 ); 
xor ( n1627 , n1281 , n1141 ); 
and ( n1628 , n1162 , n1133 ); 
not ( n1629 , n1162 ); 
and ( n1630 , n1629 , n1134 ); 
nor ( n1631 , n1628 , n1630 ); 
xnor ( n1632 , n1627 , n1631 ); 
not ( n1633 , n1632 ); 
and ( n1634 , n1171 , n1114 ); 
not ( n1635 , n1171 ); 
and ( n1636 , n1635 , n1300 ); 
or ( n1637 , n1634 , n1636 ); 
not ( n1638 , n1101 ); 
not ( n1639 , n1295 ); 
or ( n1640 , n1638 , n1639 ); 
not ( n1641 , n1101 ); 
nand ( n1642 , n1641 , n1294 ); 
nand ( n1643 , n1640 , n1642 ); 
not ( n1644 , n1125 ); 
and ( n1645 , n6 , n114 ); 
not ( n1646 , n6 ); 
and ( n1647 , n1646 , n113 ); 
nor ( n1648 , n1645 , n1647 ); 
not ( n1649 , n1648 ); 
or ( n1650 , n1644 , n1649 ); 
not ( n1651 , n1648 ); 
nand ( n1652 , n1651 , n1124 ); 
nand ( n1653 , n1650 , n1652 ); 
and ( n1654 , n1643 , n1653 ); 
not ( n1655 , n1643 ); 
not ( n1656 , n1653 ); 
and ( n1657 , n1655 , n1656 ); 
nor ( n1658 , n1654 , n1657 ); 
not ( n1659 , n1658 ); 
and ( n1660 , n1637 , n1659 ); 
not ( n1661 , n1637 ); 
and ( n1662 , n1661 , n1658 ); 
nor ( n1663 , n1660 , n1662 ); 
not ( n1664 , n1663 ); 
or ( n1665 , n1633 , n1664 ); 
or ( n1666 , n1632 , n1663 ); 
nand ( n1667 , n1665 , n1666 ); 
nand ( n1668 , n1592 , n1626 , n1667 ); 
not ( n1669 , n1668 ); 
and ( n1670 , n97 , n98 ); 
nand ( n1671 , n1670 , n96 , n99 , n100 ); 
nand ( n1672 , n102 , n103 ); 
nand ( n1673 , n101 , n104 , n105 ); 
nor ( n1674 , n1671 , n1672 , n1673 ); 
not ( n1675 , n95 ); 
and ( n1676 , n107 , n108 ); 
nand ( n1677 , n1676 , n106 , n109 , n110 ); 
not ( n1678 , n280 ); 
not ( n1679 , n235 ); 
or ( n1680 , n1678 , n1679 ); 
nand ( n1681 , n234 , n281 ); 
nand ( n1682 , n1680 , n1681 ); 
not ( n1683 , n1682 ); 
not ( n1684 , n122 ); 
and ( n1685 , n6 , n1684 ); 
not ( n1686 , n6 ); 
and ( n1687 , n1686 , n121 ); 
nor ( n1688 , n1685 , n1687 ); 
not ( n1689 , n1688 ); 
not ( n1690 , n292 ); 
and ( n1691 , n1689 , n1690 ); 
and ( n1692 , n292 , n1688 ); 
nor ( n1693 , n1691 , n1692 ); 
not ( n1694 , n1693 ); 
or ( n1695 , n1683 , n1694 ); 
or ( n1696 , n1693 , n1682 ); 
nand ( n1697 , n1695 , n1696 ); 
and ( n1698 , n308 , n262 ); 
not ( n1699 , n308 ); 
and ( n1700 , n1699 , n263 ); 
nor ( n1701 , n1698 , n1700 ); 
not ( n1702 , n1701 ); 
and ( n1703 , n1697 , n1702 ); 
not ( n1704 , n1697 ); 
and ( n1705 , n1704 , n1701 ); 
nor ( n1706 , n1703 , n1705 ); 
not ( n1707 , n4 ); 
and ( n1708 , n6 , n1707 ); 
not ( n1709 , n6 ); 
and ( n1710 , n1709 , n119 ); 
nor ( n1711 , n1708 , n1710 ); 
not ( n1712 , n1711 ); 
and ( n1713 , n6 , n2 ); 
not ( n1714 , n6 ); 
and ( n1715 , n1714 , n216 ); 
nor ( n1716 , n1713 , n1715 ); 
not ( n1717 , n1716 ); 
and ( n1718 , n1712 , n1717 ); 
and ( n1719 , n1716 , n1711 ); 
nor ( n1720 , n1718 , n1719 ); 
and ( n1721 , n1706 , n1720 ); 
not ( n1722 , n1706 ); 
not ( n1723 , n1720 ); 
and ( n1724 , n1722 , n1723 ); 
nor ( n1725 , n1721 , n1724 ); 
not ( n1726 , n567 ); 
not ( n1727 , n580 ); 
and ( n1728 , n1726 , n1727 ); 
and ( n1729 , n580 , n567 ); 
nor ( n1730 , n1728 , n1729 ); 
not ( n1731 , n1730 ); 
and ( n1732 , n553 , n536 ); 
not ( n1733 , n553 ); 
and ( n1734 , n1733 , n537 ); 
nor ( n1735 , n1732 , n1734 ); 
not ( n1736 , n1735 ); 
and ( n1737 , n1731 , n1736 ); 
and ( n1738 , n1735 , n1730 ); 
nor ( n1739 , n1737 , n1738 ); 
not ( n1740 , n483 ); 
not ( n1741 , n1740 ); 
not ( n1742 , n770 ); 
or ( n1743 , n1741 , n1742 ); 
nand ( n1744 , n769 , n483 ); 
nand ( n1745 , n1743 , n1744 ); 
not ( n1746 , n1745 ); 
not ( n1747 , n133 ); 
and ( n1748 , n6 , n1747 ); 
not ( n1749 , n6 ); 
and ( n1750 , n1749 , n132 ); 
nor ( n1751 , n1748 , n1750 ); 
not ( n1752 , n1751 ); 
not ( n1753 , n500 ); 
and ( n1754 , n1752 , n1753 ); 
and ( n1755 , n500 , n1751 ); 
nor ( n1756 , n1754 , n1755 ); 
not ( n1757 , n1756 ); 
or ( n1758 , n1746 , n1757 ); 
or ( n1759 , n1756 , n1745 ); 
nand ( n1760 , n1758 , n1759 ); 
and ( n1761 , n519 , n511 ); 
not ( n1762 , n519 ); 
and ( n1763 , n1762 , n512 ); 
or ( n1764 , n1761 , n1763 ); 
not ( n1765 , n1764 ); 
and ( n1766 , n1760 , n1765 ); 
not ( n1767 , n1760 ); 
and ( n1768 , n1767 , n1764 ); 
nor ( n1769 , n1766 , n1768 ); 
and ( n1770 , n1739 , n1769 ); 
not ( n1771 , n1739 ); 
not ( n1772 , n1769 ); 
and ( n1773 , n1771 , n1772 ); 
nor ( n1774 , n1770 , n1773 ); 
nand ( n1775 , n1725 , n1774 ); 
not ( n1776 , n335 ); 
not ( n1777 , n327 ); 
or ( n1778 , n1776 , n1777 ); 
nand ( n1779 , n325 , n334 ); 
nand ( n1780 , n1778 , n1779 ); 
and ( n1781 , n355 , n366 ); 
not ( n1782 , n355 ); 
and ( n1783 , n1782 , n367 ); 
nor ( n1784 , n1781 , n1783 ); 
xnor ( n1785 , n1780 , n1784 ); 
not ( n1786 , n1785 ); 
not ( n1787 , n798 ); 
not ( n1788 , n807 ); 
or ( n1789 , n1787 , n1788 ); 
not ( n1790 , n798 ); 
nand ( n1791 , n806 , n1790 ); 
nand ( n1792 , n1789 , n1791 ); 
and ( n1793 , n6 , n143 ); 
not ( n1794 , n6 ); 
not ( n1795 , n144 ); 
and ( n1796 , n1794 , n1795 ); 
nor ( n1797 , n1793 , n1796 ); 
not ( n1798 , n1797 ); 
not ( n1799 , n436 ); 
or ( n1800 , n1798 , n1799 ); 
or ( n1801 , n436 , n1797 ); 
nand ( n1802 , n1800 , n1801 ); 
and ( n1803 , n1792 , n1802 ); 
not ( n1804 , n1792 ); 
not ( n1805 , n1802 ); 
and ( n1806 , n1804 , n1805 ); 
nor ( n1807 , n1803 , n1806 ); 
not ( n1808 , n813 ); 
and ( n1809 , n1808 , n405 ); 
not ( n1810 , n1808 ); 
and ( n1811 , n1810 , n406 ); 
nor ( n1812 , n1809 , n1811 ); 
not ( n1813 , n1812 ); 
and ( n1814 , n1807 , n1813 ); 
not ( n1815 , n1807 ); 
and ( n1816 , n1815 , n1812 ); 
nor ( n1817 , n1814 , n1816 ); 
not ( n1818 , n1817 ); 
not ( n1819 , n1818 ); 
or ( n1820 , n1786 , n1819 ); 
not ( n1821 , n1785 ); 
nand ( n1822 , n1821 , n1817 ); 
nand ( n1823 , n1820 , n1822 ); 
not ( n1824 , n686 ); 
not ( n1825 , n652 ); 
or ( n1826 , n1824 , n1825 ); 
nand ( n1827 , n661 , n685 ); 
nand ( n1828 , n1826 , n1827 ); 
not ( n1829 , n1828 ); 
not ( n1830 , n91 ); 
nand ( n1831 , n6 , n1830 ); 
nand ( n1832 , n712 , n1831 ); 
not ( n1833 , n154 ); 
and ( n1834 , n6 , n1833 ); 
not ( n1835 , n6 ); 
and ( n1836 , n1835 , n155 ); 
nor ( n1837 , n1834 , n1836 ); 
not ( n1838 , n1837 ); 
and ( n1839 , n1832 , n1838 ); 
not ( n1840 , n1832 ); 
and ( n1841 , n1840 , n1837 ); 
nor ( n1842 , n1839 , n1841 ); 
not ( n1843 , n1842 ); 
or ( n1844 , n1829 , n1843 ); 
or ( n1845 , n1828 , n1842 ); 
nand ( n1846 , n1844 , n1845 ); 
and ( n1847 , n698 , n669 ); 
not ( n1848 , n698 ); 
and ( n1849 , n1848 , n727 ); 
nor ( n1850 , n1847 , n1849 ); 
and ( n1851 , n1846 , n1850 ); 
nor ( n1852 , n1851 , t_0 ); 
not ( n1853 , n599 ); 
not ( n1854 , n614 ); 
or ( n1855 , n1853 , n1854 ); 
nand ( n1856 , n613 , n598 ); 
nand ( n1857 , n1855 , n1856 ); 
and ( n1858 , n625 , n640 ); 
not ( n1859 , n625 ); 
and ( n1860 , n1859 , n643 ); 
nor ( n1861 , n1858 , n1860 ); 
xor ( n1862 , n1857 , n1861 ); 
not ( n1863 , n1862 ); 
and ( n1864 , n1852 , n1863 ); 
not ( n1865 , n1852 ); 
and ( n1866 , n1865 , n1862 ); 
nor ( n1867 , n1864 , n1866 ); 
nand ( n1868 , n1823 , n1867 ); 
nor ( n1869 , n1675 , n1677 , n1775 , n1868 ); 
nand ( n1870 , n1503 , n1669 , n1674 , n1869 ); 
or ( n1871 , n1775 , n1868 ); 
xor ( n1872 , n1062 , n94 ); 
not ( n1873 , n1434 ); 
patch p0 (.t_0(t_0), .g1(n684), .g2(n681), .g3(n1177), .g4(n694), .g5(n1830), .g6(n697), .g7(n712), .g8(n1201), .g9(n1833), .g10(n648), .g11(n651), .g12(n1836), .g13(n668));
endmodule 

